// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 13 2025 20:50:07

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49929;
    wire N__49928;
    wire N__49927;
    wire N__49920;
    wire N__49919;
    wire N__49918;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49902;
    wire N__49901;
    wire N__49900;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49875;
    wire N__49874;
    wire N__49873;
    wire N__49866;
    wire N__49865;
    wire N__49864;
    wire N__49857;
    wire N__49856;
    wire N__49855;
    wire N__49848;
    wire N__49847;
    wire N__49846;
    wire N__49839;
    wire N__49838;
    wire N__49837;
    wire N__49820;
    wire N__49817;
    wire N__49814;
    wire N__49811;
    wire N__49808;
    wire N__49805;
    wire N__49802;
    wire N__49799;
    wire N__49796;
    wire N__49793;
    wire N__49790;
    wire N__49787;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49779;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49772;
    wire N__49767;
    wire N__49766;
    wire N__49765;
    wire N__49764;
    wire N__49763;
    wire N__49762;
    wire N__49761;
    wire N__49758;
    wire N__49757;
    wire N__49756;
    wire N__49755;
    wire N__49754;
    wire N__49753;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49749;
    wire N__49748;
    wire N__49747;
    wire N__49746;
    wire N__49745;
    wire N__49744;
    wire N__49743;
    wire N__49742;
    wire N__49741;
    wire N__49740;
    wire N__49739;
    wire N__49738;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49733;
    wire N__49732;
    wire N__49729;
    wire N__49716;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49708;
    wire N__49707;
    wire N__49702;
    wire N__49699;
    wire N__49688;
    wire N__49685;
    wire N__49670;
    wire N__49665;
    wire N__49660;
    wire N__49655;
    wire N__49646;
    wire N__49645;
    wire N__49636;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49622;
    wire N__49621;
    wire N__49620;
    wire N__49619;
    wire N__49618;
    wire N__49617;
    wire N__49610;
    wire N__49607;
    wire N__49604;
    wire N__49599;
    wire N__49596;
    wire N__49591;
    wire N__49590;
    wire N__49589;
    wire N__49588;
    wire N__49587;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49579;
    wire N__49578;
    wire N__49577;
    wire N__49570;
    wire N__49567;
    wire N__49566;
    wire N__49565;
    wire N__49562;
    wire N__49561;
    wire N__49556;
    wire N__49539;
    wire N__49534;
    wire N__49529;
    wire N__49526;
    wire N__49523;
    wire N__49514;
    wire N__49511;
    wire N__49508;
    wire N__49499;
    wire N__49494;
    wire N__49485;
    wire N__49476;
    wire N__49457;
    wire N__49456;
    wire N__49455;
    wire N__49454;
    wire N__49451;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49443;
    wire N__49440;
    wire N__49439;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49431;
    wire N__49430;
    wire N__49429;
    wire N__49428;
    wire N__49427;
    wire N__49424;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49409;
    wire N__49406;
    wire N__49403;
    wire N__49402;
    wire N__49401;
    wire N__49400;
    wire N__49397;
    wire N__49396;
    wire N__49395;
    wire N__49394;
    wire N__49393;
    wire N__49392;
    wire N__49391;
    wire N__49390;
    wire N__49389;
    wire N__49388;
    wire N__49385;
    wire N__49382;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49377;
    wire N__49374;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49356;
    wire N__49355;
    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49351;
    wire N__49350;
    wire N__49349;
    wire N__49342;
    wire N__49337;
    wire N__49332;
    wire N__49329;
    wire N__49318;
    wire N__49315;
    wire N__49312;
    wire N__49311;
    wire N__49310;
    wire N__49309;
    wire N__49308;
    wire N__49305;
    wire N__49302;
    wire N__49299;
    wire N__49296;
    wire N__49293;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49285;
    wire N__49284;
    wire N__49283;
    wire N__49282;
    wire N__49281;
    wire N__49280;
    wire N__49279;
    wire N__49278;
    wire N__49277;
    wire N__49276;
    wire N__49275;
    wire N__49274;
    wire N__49273;
    wire N__49272;
    wire N__49267;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49256;
    wire N__49255;
    wire N__49254;
    wire N__49251;
    wire N__49250;
    wire N__49249;
    wire N__49248;
    wire N__49243;
    wire N__49236;
    wire N__49231;
    wire N__49228;
    wire N__49225;
    wire N__49224;
    wire N__49221;
    wire N__49220;
    wire N__49217;
    wire N__49216;
    wire N__49213;
    wire N__49212;
    wire N__49209;
    wire N__49208;
    wire N__49205;
    wire N__49204;
    wire N__49203;
    wire N__49202;
    wire N__49201;
    wire N__49200;
    wire N__49199;
    wire N__49198;
    wire N__49197;
    wire N__49196;
    wire N__49195;
    wire N__49192;
    wire N__49191;
    wire N__49188;
    wire N__49187;
    wire N__49184;
    wire N__49183;
    wire N__49180;
    wire N__49179;
    wire N__49178;
    wire N__49175;
    wire N__49174;
    wire N__49171;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49159;
    wire N__49154;
    wire N__49137;
    wire N__49128;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49111;
    wire N__49110;
    wire N__49107;
    wire N__49106;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49100;
    wire N__49099;
    wire N__49096;
    wire N__49095;
    wire N__49092;
    wire N__49091;
    wire N__49088;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49080;
    wire N__49077;
    wire N__49076;
    wire N__49073;
    wire N__49072;
    wire N__49069;
    wire N__49068;
    wire N__49065;
    wire N__49060;
    wire N__49055;
    wire N__49040;
    wire N__49035;
    wire N__49032;
    wire N__49021;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48995;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48984;
    wire N__48983;
    wire N__48980;
    wire N__48979;
    wire N__48976;
    wire N__48975;
    wire N__48972;
    wire N__48955;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48931;
    wire N__48926;
    wire N__48917;
    wire N__48912;
    wire N__48903;
    wire N__48900;
    wire N__48883;
    wire N__48866;
    wire N__48849;
    wire N__48840;
    wire N__48831;
    wire N__48818;
    wire N__48813;
    wire N__48782;
    wire N__48779;
    wire N__48776;
    wire N__48773;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48765;
    wire N__48760;
    wire N__48755;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48734;
    wire N__48731;
    wire N__48728;
    wire N__48725;
    wire N__48722;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48709;
    wire N__48706;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48696;
    wire N__48689;
    wire N__48688;
    wire N__48687;
    wire N__48686;
    wire N__48685;
    wire N__48680;
    wire N__48677;
    wire N__48676;
    wire N__48675;
    wire N__48674;
    wire N__48673;
    wire N__48672;
    wire N__48671;
    wire N__48670;
    wire N__48669;
    wire N__48668;
    wire N__48667;
    wire N__48666;
    wire N__48665;
    wire N__48662;
    wire N__48659;
    wire N__48658;
    wire N__48653;
    wire N__48640;
    wire N__48635;
    wire N__48630;
    wire N__48625;
    wire N__48622;
    wire N__48617;
    wire N__48614;
    wire N__48609;
    wire N__48608;
    wire N__48607;
    wire N__48606;
    wire N__48605;
    wire N__48604;
    wire N__48603;
    wire N__48598;
    wire N__48595;
    wire N__48588;
    wire N__48579;
    wire N__48576;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48559;
    wire N__48556;
    wire N__48545;
    wire N__48544;
    wire N__48541;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48531;
    wire N__48528;
    wire N__48525;
    wire N__48522;
    wire N__48519;
    wire N__48512;
    wire N__48509;
    wire N__48508;
    wire N__48505;
    wire N__48502;
    wire N__48497;
    wire N__48496;
    wire N__48495;
    wire N__48492;
    wire N__48487;
    wire N__48482;
    wire N__48481;
    wire N__48480;
    wire N__48479;
    wire N__48478;
    wire N__48477;
    wire N__48476;
    wire N__48475;
    wire N__48474;
    wire N__48473;
    wire N__48472;
    wire N__48471;
    wire N__48470;
    wire N__48469;
    wire N__48468;
    wire N__48467;
    wire N__48466;
    wire N__48465;
    wire N__48464;
    wire N__48463;
    wire N__48462;
    wire N__48461;
    wire N__48460;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48456;
    wire N__48455;
    wire N__48454;
    wire N__48453;
    wire N__48452;
    wire N__48451;
    wire N__48450;
    wire N__48449;
    wire N__48448;
    wire N__48447;
    wire N__48446;
    wire N__48445;
    wire N__48444;
    wire N__48443;
    wire N__48442;
    wire N__48441;
    wire N__48440;
    wire N__48439;
    wire N__48438;
    wire N__48437;
    wire N__48436;
    wire N__48435;
    wire N__48434;
    wire N__48433;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48426;
    wire N__48425;
    wire N__48424;
    wire N__48423;
    wire N__48422;
    wire N__48421;
    wire N__48420;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48399;
    wire N__48398;
    wire N__48397;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48390;
    wire N__48389;
    wire N__48388;
    wire N__48387;
    wire N__48386;
    wire N__48385;
    wire N__48384;
    wire N__48383;
    wire N__48382;
    wire N__48381;
    wire N__48380;
    wire N__48379;
    wire N__48378;
    wire N__48377;
    wire N__48376;
    wire N__48375;
    wire N__48374;
    wire N__48373;
    wire N__48372;
    wire N__48371;
    wire N__48370;
    wire N__48369;
    wire N__48368;
    wire N__48367;
    wire N__48366;
    wire N__48365;
    wire N__48364;
    wire N__48363;
    wire N__48362;
    wire N__48361;
    wire N__48360;
    wire N__48359;
    wire N__48358;
    wire N__48357;
    wire N__48356;
    wire N__48355;
    wire N__48354;
    wire N__48353;
    wire N__48352;
    wire N__48351;
    wire N__48350;
    wire N__48349;
    wire N__48348;
    wire N__48347;
    wire N__48346;
    wire N__48345;
    wire N__48344;
    wire N__48343;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48336;
    wire N__48335;
    wire N__48334;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48330;
    wire N__48329;
    wire N__48020;
    wire N__48017;
    wire N__48016;
    wire N__48013;
    wire N__48012;
    wire N__48009;
    wire N__48008;
    wire N__48005;
    wire N__48002;
    wire N__47999;
    wire N__47996;
    wire N__47995;
    wire N__47994;
    wire N__47989;
    wire N__47988;
    wire N__47987;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47960;
    wire N__47955;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47942;
    wire N__47937;
    wire N__47932;
    wire N__47927;
    wire N__47926;
    wire N__47925;
    wire N__47924;
    wire N__47923;
    wire N__47922;
    wire N__47919;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47885;
    wire N__47884;
    wire N__47883;
    wire N__47882;
    wire N__47881;
    wire N__47880;
    wire N__47879;
    wire N__47878;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47860;
    wire N__47859;
    wire N__47858;
    wire N__47857;
    wire N__47856;
    wire N__47855;
    wire N__47854;
    wire N__47853;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47844;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47830;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47826;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47812;
    wire N__47811;
    wire N__47810;
    wire N__47809;
    wire N__47808;
    wire N__47807;
    wire N__47806;
    wire N__47805;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47801;
    wire N__47800;
    wire N__47799;
    wire N__47798;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47790;
    wire N__47789;
    wire N__47788;
    wire N__47787;
    wire N__47786;
    wire N__47785;
    wire N__47784;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47776;
    wire N__47775;
    wire N__47774;
    wire N__47773;
    wire N__47772;
    wire N__47771;
    wire N__47770;
    wire N__47769;
    wire N__47768;
    wire N__47767;
    wire N__47766;
    wire N__47765;
    wire N__47762;
    wire N__47761;
    wire N__47760;
    wire N__47759;
    wire N__47758;
    wire N__47757;
    wire N__47756;
    wire N__47755;
    wire N__47754;
    wire N__47753;
    wire N__47752;
    wire N__47751;
    wire N__47750;
    wire N__47749;
    wire N__47748;
    wire N__47747;
    wire N__47746;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47740;
    wire N__47739;
    wire N__47738;
    wire N__47737;
    wire N__47736;
    wire N__47735;
    wire N__47444;
    wire N__47441;
    wire N__47438;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47427;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47417;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47403;
    wire N__47398;
    wire N__47395;
    wire N__47390;
    wire N__47387;
    wire N__47386;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47376;
    wire N__47369;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47336;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47318;
    wire N__47317;
    wire N__47314;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47297;
    wire N__47294;
    wire N__47291;
    wire N__47288;
    wire N__47287;
    wire N__47286;
    wire N__47283;
    wire N__47282;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47260;
    wire N__47255;
    wire N__47254;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47237;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47227;
    wire N__47224;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47206;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47189;
    wire N__47186;
    wire N__47185;
    wire N__47184;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47168;
    wire N__47165;
    wire N__47162;
    wire N__47159;
    wire N__47158;
    wire N__47155;
    wire N__47152;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47137;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47116;
    wire N__47115;
    wire N__47110;
    wire N__47107;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47095;
    wire N__47094;
    wire N__47091;
    wire N__47088;
    wire N__47085;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47068;
    wire N__47067;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47054;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47037;
    wire N__47034;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47008;
    wire N__47005;
    wire N__47004;
    wire N__47001;
    wire N__46996;
    wire N__46991;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46979;
    wire N__46978;
    wire N__46977;
    wire N__46974;
    wire N__46969;
    wire N__46964;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46956;
    wire N__46951;
    wire N__46948;
    wire N__46945;
    wire N__46942;
    wire N__46937;
    wire N__46934;
    wire N__46931;
    wire N__46930;
    wire N__46927;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46905;
    wire N__46904;
    wire N__46901;
    wire N__46896;
    wire N__46893;
    wire N__46886;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46865;
    wire N__46862;
    wire N__46859;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46832;
    wire N__46829;
    wire N__46824;
    wire N__46821;
    wire N__46814;
    wire N__46811;
    wire N__46810;
    wire N__46809;
    wire N__46806;
    wire N__46803;
    wire N__46800;
    wire N__46793;
    wire N__46790;
    wire N__46787;
    wire N__46784;
    wire N__46783;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46754;
    wire N__46751;
    wire N__46746;
    wire N__46743;
    wire N__46736;
    wire N__46733;
    wire N__46732;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46702;
    wire N__46701;
    wire N__46698;
    wire N__46695;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46685;
    wire N__46682;
    wire N__46679;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46667;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46649;
    wire N__46648;
    wire N__46645;
    wire N__46642;
    wire N__46639;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46622;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46612;
    wire N__46611;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46593;
    wire N__46588;
    wire N__46585;
    wire N__46580;
    wire N__46579;
    wire N__46578;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46562;
    wire N__46559;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46546;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46530;
    wire N__46527;
    wire N__46522;
    wire N__46521;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46505;
    wire N__46502;
    wire N__46501;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46475;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46462;
    wire N__46461;
    wire N__46460;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46446;
    wire N__46445;
    wire N__46444;
    wire N__46443;
    wire N__46442;
    wire N__46441;
    wire N__46440;
    wire N__46439;
    wire N__46438;
    wire N__46433;
    wire N__46430;
    wire N__46413;
    wire N__46406;
    wire N__46403;
    wire N__46400;
    wire N__46397;
    wire N__46394;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46366;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46354;
    wire N__46353;
    wire N__46350;
    wire N__46349;
    wire N__46346;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46310;
    wire N__46307;
    wire N__46304;
    wire N__46303;
    wire N__46302;
    wire N__46295;
    wire N__46292;
    wire N__46291;
    wire N__46290;
    wire N__46289;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46268;
    wire N__46267;
    wire N__46266;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46238;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46220;
    wire N__46219;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46192;
    wire N__46187;
    wire N__46184;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46151;
    wire N__46150;
    wire N__46149;
    wire N__46148;
    wire N__46147;
    wire N__46146;
    wire N__46145;
    wire N__46142;
    wire N__46139;
    wire N__46136;
    wire N__46133;
    wire N__46130;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46122;
    wire N__46121;
    wire N__46120;
    wire N__46119;
    wire N__46118;
    wire N__46117;
    wire N__46116;
    wire N__46115;
    wire N__46114;
    wire N__46113;
    wire N__46104;
    wire N__46095;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46042;
    wire N__46041;
    wire N__46040;
    wire N__46039;
    wire N__46038;
    wire N__46037;
    wire N__46036;
    wire N__46035;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46028;
    wire N__46027;
    wire N__46026;
    wire N__46025;
    wire N__46024;
    wire N__46017;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45983;
    wire N__45980;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45967;
    wire N__45966;
    wire N__45963;
    wire N__45956;
    wire N__45947;
    wire N__45942;
    wire N__45935;
    wire N__45932;
    wire N__45925;
    wire N__45916;
    wire N__45913;
    wire N__45912;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45904;
    wire N__45897;
    wire N__45896;
    wire N__45895;
    wire N__45894;
    wire N__45893;
    wire N__45892;
    wire N__45891;
    wire N__45890;
    wire N__45889;
    wire N__45878;
    wire N__45875;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45861;
    wire N__45858;
    wire N__45857;
    wire N__45856;
    wire N__45849;
    wire N__45840;
    wire N__45837;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45805;
    wire N__45800;
    wire N__45795;
    wire N__45790;
    wire N__45787;
    wire N__45782;
    wire N__45779;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45759;
    wire N__45752;
    wire N__45749;
    wire N__45746;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45728;
    wire N__45725;
    wire N__45722;
    wire N__45719;
    wire N__45716;
    wire N__45713;
    wire N__45710;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45667;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45657;
    wire N__45650;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45617;
    wire N__45616;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45599;
    wire N__45596;
    wire N__45595;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45580;
    wire N__45577;
    wire N__45574;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45566;
    wire N__45565;
    wire N__45564;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45496;
    wire N__45493;
    wire N__45488;
    wire N__45487;
    wire N__45486;
    wire N__45483;
    wire N__45482;
    wire N__45481;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45459;
    wire N__45458;
    wire N__45455;
    wire N__45452;
    wire N__45449;
    wire N__45446;
    wire N__45439;
    wire N__45434;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45404;
    wire N__45401;
    wire N__45398;
    wire N__45397;
    wire N__45396;
    wire N__45393;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45368;
    wire N__45365;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45326;
    wire N__45325;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45295;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45283;
    wire N__45282;
    wire N__45281;
    wire N__45278;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45232;
    wire N__45231;
    wire N__45228;
    wire N__45227;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45172;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45154;
    wire N__45149;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45137;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45115;
    wire N__45114;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45068;
    wire N__45065;
    wire N__45062;
    wire N__45059;
    wire N__45056;
    wire N__45053;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45023;
    wire N__45020;
    wire N__45019;
    wire N__45018;
    wire N__45015;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44977;
    wire N__44976;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44960;
    wire N__44957;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44906;
    wire N__44903;
    wire N__44902;
    wire N__44899;
    wire N__44898;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44882;
    wire N__44879;
    wire N__44876;
    wire N__44873;
    wire N__44870;
    wire N__44867;
    wire N__44864;
    wire N__44861;
    wire N__44858;
    wire N__44855;
    wire N__44852;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44825;
    wire N__44822;
    wire N__44821;
    wire N__44818;
    wire N__44817;
    wire N__44814;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44798;
    wire N__44795;
    wire N__44794;
    wire N__44789;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44762;
    wire N__44759;
    wire N__44758;
    wire N__44757;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44741;
    wire N__44738;
    wire N__44737;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44717;
    wire N__44714;
    wire N__44711;
    wire N__44708;
    wire N__44705;
    wire N__44704;
    wire N__44703;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44678;
    wire N__44675;
    wire N__44672;
    wire N__44671;
    wire N__44668;
    wire N__44665;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44647;
    wire N__44642;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44630;
    wire N__44627;
    wire N__44626;
    wire N__44623;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44572;
    wire N__44571;
    wire N__44568;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44540;
    wire N__44537;
    wire N__44536;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44508;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44461;
    wire N__44460;
    wire N__44457;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44416;
    wire N__44413;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44396;
    wire N__44393;
    wire N__44388;
    wire N__44385;
    wire N__44378;
    wire N__44377;
    wire N__44376;
    wire N__44373;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44339;
    wire N__44336;
    wire N__44335;
    wire N__44334;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44318;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44263;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44237;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44167;
    wire N__44162;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44151;
    wire N__44146;
    wire N__44143;
    wire N__44138;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44119;
    wire N__44118;
    wire N__44117;
    wire N__44116;
    wire N__44115;
    wire N__44114;
    wire N__44113;
    wire N__44104;
    wire N__44095;
    wire N__44094;
    wire N__44093;
    wire N__44092;
    wire N__44091;
    wire N__44090;
    wire N__44089;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44085;
    wire N__44084;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44077;
    wire N__44072;
    wire N__44063;
    wire N__44058;
    wire N__44057;
    wire N__44056;
    wire N__44055;
    wire N__44054;
    wire N__44045;
    wire N__44036;
    wire N__44027;
    wire N__44020;
    wire N__44011;
    wire N__44006;
    wire N__44001;
    wire N__43998;
    wire N__43993;
    wire N__43988;
    wire N__43985;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43973;
    wire N__43970;
    wire N__43969;
    wire N__43966;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43955;
    wire N__43948;
    wire N__43945;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43916;
    wire N__43915;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43900;
    wire N__43895;
    wire N__43892;
    wire N__43889;
    wire N__43886;
    wire N__43883;
    wire N__43882;
    wire N__43881;
    wire N__43880;
    wire N__43879;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43863;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43826;
    wire N__43825;
    wire N__43824;
    wire N__43823;
    wire N__43822;
    wire N__43821;
    wire N__43820;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43816;
    wire N__43815;
    wire N__43808;
    wire N__43805;
    wire N__43804;
    wire N__43801;
    wire N__43800;
    wire N__43799;
    wire N__43798;
    wire N__43797;
    wire N__43796;
    wire N__43795;
    wire N__43794;
    wire N__43779;
    wire N__43778;
    wire N__43777;
    wire N__43776;
    wire N__43775;
    wire N__43772;
    wire N__43767;
    wire N__43750;
    wire N__43747;
    wire N__43738;
    wire N__43735;
    wire N__43724;
    wire N__43723;
    wire N__43722;
    wire N__43721;
    wire N__43720;
    wire N__43719;
    wire N__43718;
    wire N__43717;
    wire N__43716;
    wire N__43713;
    wire N__43712;
    wire N__43709;
    wire N__43708;
    wire N__43705;
    wire N__43704;
    wire N__43701;
    wire N__43700;
    wire N__43697;
    wire N__43696;
    wire N__43695;
    wire N__43692;
    wire N__43691;
    wire N__43688;
    wire N__43687;
    wire N__43684;
    wire N__43683;
    wire N__43678;
    wire N__43661;
    wire N__43660;
    wire N__43657;
    wire N__43644;
    wire N__43641;
    wire N__43640;
    wire N__43635;
    wire N__43634;
    wire N__43631;
    wire N__43630;
    wire N__43629;
    wire N__43624;
    wire N__43619;
    wire N__43616;
    wire N__43607;
    wire N__43602;
    wire N__43601;
    wire N__43596;
    wire N__43593;
    wire N__43590;
    wire N__43587;
    wire N__43584;
    wire N__43577;
    wire N__43576;
    wire N__43575;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43565;
    wire N__43564;
    wire N__43563;
    wire N__43562;
    wire N__43561;
    wire N__43560;
    wire N__43559;
    wire N__43558;
    wire N__43557;
    wire N__43556;
    wire N__43555;
    wire N__43554;
    wire N__43547;
    wire N__43538;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43519;
    wire N__43518;
    wire N__43517;
    wire N__43516;
    wire N__43515;
    wire N__43514;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43506;
    wire N__43497;
    wire N__43488;
    wire N__43483;
    wire N__43480;
    wire N__43471;
    wire N__43464;
    wire N__43461;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43403;
    wire N__43402;
    wire N__43401;
    wire N__43398;
    wire N__43393;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43381;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43334;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43322;
    wire N__43321;
    wire N__43320;
    wire N__43317;
    wire N__43312;
    wire N__43307;
    wire N__43304;
    wire N__43303;
    wire N__43302;
    wire N__43299;
    wire N__43294;
    wire N__43289;
    wire N__43286;
    wire N__43285;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43270;
    wire N__43265;
    wire N__43262;
    wire N__43261;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43246;
    wire N__43241;
    wire N__43238;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43217;
    wire N__43214;
    wire N__43213;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43193;
    wire N__43190;
    wire N__43189;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43174;
    wire N__43169;
    wire N__43166;
    wire N__43165;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43155;
    wire N__43150;
    wire N__43145;
    wire N__43142;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43130;
    wire N__43127;
    wire N__43126;
    wire N__43125;
    wire N__43122;
    wire N__43117;
    wire N__43112;
    wire N__43109;
    wire N__43108;
    wire N__43107;
    wire N__43104;
    wire N__43099;
    wire N__43094;
    wire N__43091;
    wire N__43090;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43075;
    wire N__43070;
    wire N__43067;
    wire N__43066;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43051;
    wire N__43046;
    wire N__43043;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43022;
    wire N__43019;
    wire N__43018;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__42998;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42979;
    wire N__42974;
    wire N__42971;
    wire N__42970;
    wire N__42969;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42955;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42943;
    wire N__42942;
    wire N__42939;
    wire N__42934;
    wire N__42929;
    wire N__42926;
    wire N__42925;
    wire N__42924;
    wire N__42921;
    wire N__42916;
    wire N__42911;
    wire N__42908;
    wire N__42907;
    wire N__42906;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42892;
    wire N__42887;
    wire N__42884;
    wire N__42883;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42868;
    wire N__42863;
    wire N__42860;
    wire N__42859;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42839;
    wire N__42836;
    wire N__42835;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42815;
    wire N__42812;
    wire N__42811;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42796;
    wire N__42791;
    wire N__42788;
    wire N__42787;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42772;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42747;
    wire N__42746;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42709;
    wire N__42706;
    wire N__42705;
    wire N__42702;
    wire N__42701;
    wire N__42700;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42687;
    wire N__42684;
    wire N__42683;
    wire N__42680;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42625;
    wire N__42620;
    wire N__42617;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42590;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42582;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42544;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42529;
    wire N__42524;
    wire N__42521;
    wire N__42520;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42505;
    wire N__42500;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42492;
    wire N__42489;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42395;
    wire N__42392;
    wire N__42389;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42338;
    wire N__42335;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42254;
    wire N__42251;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42170;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42110;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42098;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42088;
    wire N__42085;
    wire N__42082;
    wire N__42077;
    wire N__42074;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42064;
    wire N__42061;
    wire N__42058;
    wire N__42055;
    wire N__42052;
    wire N__42049;
    wire N__42044;
    wire N__42043;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42019;
    wire N__42014;
    wire N__42011;
    wire N__42008;
    wire N__42005;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41966;
    wire N__41963;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41953;
    wire N__41950;
    wire N__41947;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41933;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41909;
    wire N__41906;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41884;
    wire N__41881;
    wire N__41876;
    wire N__41873;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41759;
    wire N__41756;
    wire N__41753;
    wire N__41750;
    wire N__41747;
    wire N__41744;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41726;
    wire N__41723;
    wire N__41720;
    wire N__41717;
    wire N__41714;
    wire N__41713;
    wire N__41710;
    wire N__41707;
    wire N__41704;
    wire N__41701;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41666;
    wire N__41663;
    wire N__41660;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41650;
    wire N__41647;
    wire N__41644;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41483;
    wire N__41480;
    wire N__41477;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41434;
    wire N__41433;
    wire N__41430;
    wire N__41429;
    wire N__41428;
    wire N__41427;
    wire N__41418;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41410;
    wire N__41409;
    wire N__41408;
    wire N__41407;
    wire N__41406;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41383;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41371;
    wire N__41368;
    wire N__41365;
    wire N__41360;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41319;
    wire N__41314;
    wire N__41311;
    wire N__41306;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41281;
    wire N__41280;
    wire N__41277;
    wire N__41272;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41258;
    wire N__41257;
    wire N__41256;
    wire N__41253;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41237;
    wire N__41234;
    wire N__41233;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41132;
    wire N__41129;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41121;
    wire N__41116;
    wire N__41113;
    wire N__41112;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41088;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41057;
    wire N__41054;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41042;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40984;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40976;
    wire N__40975;
    wire N__40972;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40940;
    wire N__40937;
    wire N__40936;
    wire N__40935;
    wire N__40934;
    wire N__40929;
    wire N__40928;
    wire N__40925;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40896;
    wire N__40893;
    wire N__40888;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40873;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40834;
    wire N__40833;
    wire N__40830;
    wire N__40829;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40800;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40775;
    wire N__40772;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40730;
    wire N__40727;
    wire N__40724;
    wire N__40721;
    wire N__40718;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40706;
    wire N__40703;
    wire N__40702;
    wire N__40701;
    wire N__40700;
    wire N__40697;
    wire N__40696;
    wire N__40693;
    wire N__40692;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40680;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40661;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40640;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40613;
    wire N__40610;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40598;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40583;
    wire N__40580;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40572;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40556;
    wire N__40553;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40545;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40529;
    wire N__40526;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40518;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40502;
    wire N__40499;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40487;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40472;
    wire N__40469;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40457;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40426;
    wire N__40421;
    wire N__40418;
    wire N__40417;
    wire N__40416;
    wire N__40415;
    wire N__40414;
    wire N__40413;
    wire N__40412;
    wire N__40411;
    wire N__40410;
    wire N__40409;
    wire N__40408;
    wire N__40407;
    wire N__40406;
    wire N__40405;
    wire N__40404;
    wire N__40403;
    wire N__40402;
    wire N__40401;
    wire N__40396;
    wire N__40387;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40383;
    wire N__40382;
    wire N__40381;
    wire N__40380;
    wire N__40379;
    wire N__40378;
    wire N__40377;
    wire N__40376;
    wire N__40375;
    wire N__40366;
    wire N__40357;
    wire N__40348;
    wire N__40343;
    wire N__40334;
    wire N__40325;
    wire N__40316;
    wire N__40307;
    wire N__40298;
    wire N__40295;
    wire N__40292;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40277;
    wire N__40276;
    wire N__40275;
    wire N__40274;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40251;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40235;
    wire N__40232;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40220;
    wire N__40219;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40205;
    wire N__40202;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40194;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40178;
    wire N__40175;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40153;
    wire N__40148;
    wire N__40145;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40133;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40118;
    wire N__40115;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40103;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40088;
    wire N__40085;
    wire N__40084;
    wire N__40083;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40067;
    wire N__40064;
    wire N__40063;
    wire N__40058;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40043;
    wire N__40040;
    wire N__40039;
    wire N__40034;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40019;
    wire N__40016;
    wire N__40015;
    wire N__40010;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39995;
    wire N__39992;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39981;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39965;
    wire N__39962;
    wire N__39961;
    wire N__39958;
    wire N__39955;
    wire N__39952;
    wire N__39951;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39935;
    wire N__39932;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39920;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39905;
    wire N__39902;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39894;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39878;
    wire N__39875;
    wire N__39874;
    wire N__39873;
    wire N__39868;
    wire N__39865;
    wire N__39862;
    wire N__39857;
    wire N__39854;
    wire N__39853;
    wire N__39852;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39817;
    wire N__39816;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39800;
    wire N__39797;
    wire N__39796;
    wire N__39791;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39781;
    wire N__39776;
    wire N__39773;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39765;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39749;
    wire N__39746;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39738;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39644;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39464;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39359;
    wire N__39356;
    wire N__39353;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39332;
    wire N__39331;
    wire N__39328;
    wire N__39327;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39297;
    wire N__39294;
    wire N__39287;
    wire N__39286;
    wire N__39281;
    wire N__39278;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39260;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39252;
    wire N__39251;
    wire N__39250;
    wire N__39249;
    wire N__39248;
    wire N__39247;
    wire N__39244;
    wire N__39237;
    wire N__39232;
    wire N__39227;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39206;
    wire N__39205;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39190;
    wire N__39189;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39114;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39072;
    wire N__39067;
    wire N__39064;
    wire N__39063;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39037;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38810;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38798;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38749;
    wire N__38748;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38717;
    wire N__38714;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38706;
    wire N__38701;
    wire N__38698;
    wire N__38693;
    wire N__38692;
    wire N__38689;
    wire N__38688;
    wire N__38687;
    wire N__38686;
    wire N__38683;
    wire N__38680;
    wire N__38677;
    wire N__38672;
    wire N__38669;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38645;
    wire N__38644;
    wire N__38643;
    wire N__38642;
    wire N__38641;
    wire N__38636;
    wire N__38631;
    wire N__38628;
    wire N__38627;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38613;
    wire N__38612;
    wire N__38611;
    wire N__38608;
    wire N__38603;
    wire N__38598;
    wire N__38591;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38558;
    wire N__38557;
    wire N__38552;
    wire N__38551;
    wire N__38550;
    wire N__38549;
    wire N__38546;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38516;
    wire N__38513;
    wire N__38506;
    wire N__38501;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38492;
    wire N__38489;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38472;
    wire N__38471;
    wire N__38468;
    wire N__38463;
    wire N__38462;
    wire N__38457;
    wire N__38454;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38436;
    wire N__38431;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38393;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38375;
    wire N__38372;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38360;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38314;
    wire N__38313;
    wire N__38312;
    wire N__38311;
    wire N__38308;
    wire N__38307;
    wire N__38298;
    wire N__38297;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38285;
    wire N__38282;
    wire N__38277;
    wire N__38276;
    wire N__38275;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38258;
    wire N__38249;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38241;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38210;
    wire N__38209;
    wire N__38208;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38186;
    wire N__38183;
    wire N__38182;
    wire N__38181;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38173;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38102;
    wire N__38101;
    wire N__38100;
    wire N__38099;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38088;
    wire N__38081;
    wire N__38078;
    wire N__38069;
    wire N__38068;
    wire N__38067;
    wire N__38060;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38046;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38032;
    wire N__38027;
    wire N__38022;
    wire N__38019;
    wire N__38014;
    wire N__38009;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37997;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37989;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37834;
    wire N__37831;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37814;
    wire N__37813;
    wire N__37812;
    wire N__37811;
    wire N__37810;
    wire N__37809;
    wire N__37806;
    wire N__37805;
    wire N__37804;
    wire N__37803;
    wire N__37802;
    wire N__37801;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37793;
    wire N__37792;
    wire N__37791;
    wire N__37790;
    wire N__37789;
    wire N__37788;
    wire N__37787;
    wire N__37786;
    wire N__37785;
    wire N__37784;
    wire N__37783;
    wire N__37776;
    wire N__37773;
    wire N__37760;
    wire N__37755;
    wire N__37746;
    wire N__37739;
    wire N__37734;
    wire N__37731;
    wire N__37730;
    wire N__37727;
    wire N__37722;
    wire N__37719;
    wire N__37710;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37694;
    wire N__37685;
    wire N__37684;
    wire N__37683;
    wire N__37682;
    wire N__37681;
    wire N__37678;
    wire N__37677;
    wire N__37676;
    wire N__37675;
    wire N__37674;
    wire N__37673;
    wire N__37672;
    wire N__37671;
    wire N__37668;
    wire N__37667;
    wire N__37666;
    wire N__37665;
    wire N__37656;
    wire N__37653;
    wire N__37652;
    wire N__37651;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37631;
    wire N__37630;
    wire N__37623;
    wire N__37622;
    wire N__37619;
    wire N__37618;
    wire N__37613;
    wire N__37600;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37582;
    wire N__37577;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37538;
    wire N__37529;
    wire N__37528;
    wire N__37527;
    wire N__37526;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37522;
    wire N__37519;
    wire N__37518;
    wire N__37517;
    wire N__37516;
    wire N__37515;
    wire N__37514;
    wire N__37513;
    wire N__37512;
    wire N__37511;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37493;
    wire N__37492;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37483;
    wire N__37470;
    wire N__37467;
    wire N__37462;
    wire N__37457;
    wire N__37454;
    wire N__37445;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37437;
    wire N__37432;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37403;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37370;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37276;
    wire N__37275;
    wire N__37274;
    wire N__37273;
    wire N__37266;
    wire N__37263;
    wire N__37262;
    wire N__37261;
    wire N__37258;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37246;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37232;
    wire N__37229;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37169;
    wire N__37166;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37003;
    wire N__37002;
    wire N__37001;
    wire N__36998;
    wire N__36993;
    wire N__36990;
    wire N__36983;
    wire N__36982;
    wire N__36981;
    wire N__36980;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36917;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36861;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36850;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36808;
    wire N__36807;
    wire N__36806;
    wire N__36803;
    wire N__36798;
    wire N__36795;
    wire N__36790;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36628;
    wire N__36627;
    wire N__36626;
    wire N__36623;
    wire N__36622;
    wire N__36621;
    wire N__36620;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36604;
    wire N__36603;
    wire N__36602;
    wire N__36601;
    wire N__36598;
    wire N__36583;
    wire N__36580;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36552;
    wire N__36551;
    wire N__36550;
    wire N__36549;
    wire N__36544;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36510;
    wire N__36505;
    wire N__36502;
    wire N__36493;
    wire N__36482;
    wire N__36481;
    wire N__36480;
    wire N__36479;
    wire N__36478;
    wire N__36477;
    wire N__36476;
    wire N__36475;
    wire N__36474;
    wire N__36473;
    wire N__36472;
    wire N__36471;
    wire N__36470;
    wire N__36469;
    wire N__36468;
    wire N__36467;
    wire N__36466;
    wire N__36465;
    wire N__36464;
    wire N__36463;
    wire N__36460;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36431;
    wire N__36428;
    wire N__36427;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36380;
    wire N__36377;
    wire N__36376;
    wire N__36373;
    wire N__36366;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36332;
    wire N__36331;
    wire N__36330;
    wire N__36329;
    wire N__36328;
    wire N__36327;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36318;
    wire N__36317;
    wire N__36316;
    wire N__36315;
    wire N__36312;
    wire N__36297;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36289;
    wire N__36288;
    wire N__36287;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36254;
    wire N__36253;
    wire N__36250;
    wire N__36245;
    wire N__36238;
    wire N__36235;
    wire N__36230;
    wire N__36225;
    wire N__36212;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36164;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36148;
    wire N__36147;
    wire N__36144;
    wire N__36141;
    wire N__36138;
    wire N__36131;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36123;
    wire N__36122;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36076;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36039;
    wire N__36036;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35913;
    wire N__35908;
    wire N__35905;
    wire N__35904;
    wire N__35901;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35823;
    wire N__35822;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35810;
    wire N__35805;
    wire N__35802;
    wire N__35799;
    wire N__35796;
    wire N__35789;
    wire N__35786;
    wire N__35785;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35745;
    wire N__35742;
    wire N__35737;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35683;
    wire N__35680;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35609;
    wire N__35602;
    wire N__35601;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35585;
    wire N__35584;
    wire N__35583;
    wire N__35582;
    wire N__35581;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35575;
    wire N__35574;
    wire N__35573;
    wire N__35572;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35549;
    wire N__35548;
    wire N__35547;
    wire N__35546;
    wire N__35545;
    wire N__35544;
    wire N__35543;
    wire N__35542;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35527;
    wire N__35520;
    wire N__35503;
    wire N__35502;
    wire N__35493;
    wire N__35492;
    wire N__35491;
    wire N__35488;
    wire N__35479;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35463;
    wire N__35460;
    wire N__35455;
    wire N__35450;
    wire N__35441;
    wire N__35440;
    wire N__35439;
    wire N__35438;
    wire N__35437;
    wire N__35436;
    wire N__35435;
    wire N__35434;
    wire N__35433;
    wire N__35432;
    wire N__35431;
    wire N__35430;
    wire N__35429;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35425;
    wire N__35424;
    wire N__35423;
    wire N__35422;
    wire N__35407;
    wire N__35390;
    wire N__35381;
    wire N__35378;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35355;
    wire N__35352;
    wire N__35345;
    wire N__35340;
    wire N__35335;
    wire N__35330;
    wire N__35329;
    wire N__35328;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35291;
    wire N__35290;
    wire N__35289;
    wire N__35288;
    wire N__35279;
    wire N__35270;
    wire N__35255;
    wire N__35250;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35229;
    wire N__35226;
    wire N__35223;
    wire N__35216;
    wire N__35215;
    wire N__35214;
    wire N__35211;
    wire N__35206;
    wire N__35203;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35170;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35144;
    wire N__35141;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35133;
    wire N__35128;
    wire N__35125;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35096;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35069;
    wire N__35066;
    wire N__35065;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35039;
    wire N__35038;
    wire N__35037;
    wire N__35034;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35016;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34982;
    wire N__34979;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34971;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34952;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34940;
    wire N__34939;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34864;
    wire N__34861;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34608;
    wire N__34603;
    wire N__34600;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34560;
    wire N__34557;
    wire N__34552;
    wire N__34547;
    wire N__34546;
    wire N__34545;
    wire N__34544;
    wire N__34537;
    wire N__34534;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34503;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34425;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34401;
    wire N__34400;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34363;
    wire N__34362;
    wire N__34361;
    wire N__34360;
    wire N__34359;
    wire N__34358;
    wire N__34357;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34343;
    wire N__34342;
    wire N__34341;
    wire N__34340;
    wire N__34339;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34329;
    wire N__34326;
    wire N__34309;
    wire N__34304;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34295;
    wire N__34294;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34290;
    wire N__34289;
    wire N__34288;
    wire N__34285;
    wire N__34284;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34268;
    wire N__34267;
    wire N__34266;
    wire N__34265;
    wire N__34264;
    wire N__34259;
    wire N__34250;
    wire N__34239;
    wire N__34234;
    wire N__34227;
    wire N__34224;
    wire N__34211;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34184;
    wire N__34183;
    wire N__34178;
    wire N__34177;
    wire N__34176;
    wire N__34175;
    wire N__34174;
    wire N__34173;
    wire N__34172;
    wire N__34171;
    wire N__34170;
    wire N__34169;
    wire N__34168;
    wire N__34167;
    wire N__34166;
    wire N__34165;
    wire N__34162;
    wire N__34157;
    wire N__34156;
    wire N__34155;
    wire N__34142;
    wire N__34131;
    wire N__34130;
    wire N__34129;
    wire N__34128;
    wire N__34123;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34105;
    wire N__34104;
    wire N__34103;
    wire N__34102;
    wire N__34101;
    wire N__34100;
    wire N__34099;
    wire N__34098;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34084;
    wire N__34067;
    wire N__34058;
    wire N__34055;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34044;
    wire N__34043;
    wire N__34040;
    wire N__34039;
    wire N__34036;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34020;
    wire N__34013;
    wire N__34012;
    wire N__34011;
    wire N__34010;
    wire N__34009;
    wire N__34008;
    wire N__34005;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33992;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33976;
    wire N__33967;
    wire N__33964;
    wire N__33963;
    wire N__33962;
    wire N__33961;
    wire N__33960;
    wire N__33959;
    wire N__33958;
    wire N__33957;
    wire N__33956;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33948;
    wire N__33947;
    wire N__33946;
    wire N__33945;
    wire N__33942;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33928;
    wire N__33927;
    wire N__33924;
    wire N__33923;
    wire N__33922;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33911;
    wire N__33910;
    wire N__33909;
    wire N__33908;
    wire N__33907;
    wire N__33904;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33867;
    wire N__33858;
    wire N__33841;
    wire N__33836;
    wire N__33831;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33799;
    wire N__33798;
    wire N__33795;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33773;
    wire N__33770;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33751;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33743;
    wire N__33740;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33728;
    wire N__33725;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33704;
    wire N__33703;
    wire N__33702;
    wire N__33699;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33654;
    wire N__33651;
    wire N__33644;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33619;
    wire N__33616;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33598;
    wire N__33593;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33585;
    wire N__33582;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33548;
    wire N__33545;
    wire N__33540;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33520;
    wire N__33519;
    wire N__33518;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33514;
    wire N__33513;
    wire N__33512;
    wire N__33511;
    wire N__33510;
    wire N__33509;
    wire N__33508;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33500;
    wire N__33499;
    wire N__33496;
    wire N__33491;
    wire N__33482;
    wire N__33479;
    wire N__33478;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33474;
    wire N__33473;
    wire N__33470;
    wire N__33465;
    wire N__33460;
    wire N__33453;
    wire N__33452;
    wire N__33451;
    wire N__33448;
    wire N__33443;
    wire N__33438;
    wire N__33437;
    wire N__33432;
    wire N__33429;
    wire N__33418;
    wire N__33415;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33397;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33359;
    wire N__33354;
    wire N__33349;
    wire N__33344;
    wire N__33341;
    wire N__33326;
    wire N__33325;
    wire N__33324;
    wire N__33323;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33312;
    wire N__33309;
    wire N__33308;
    wire N__33307;
    wire N__33302;
    wire N__33297;
    wire N__33294;
    wire N__33293;
    wire N__33290;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33268;
    wire N__33263;
    wire N__33262;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33252;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33231;
    wire N__33224;
    wire N__33217;
    wire N__33212;
    wire N__33207;
    wire N__33206;
    wire N__33205;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33197;
    wire N__33188;
    wire N__33185;
    wire N__33180;
    wire N__33177;
    wire N__33172;
    wire N__33163;
    wire N__33160;
    wire N__33143;
    wire N__33142;
    wire N__33141;
    wire N__33140;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33133;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33124;
    wire N__33123;
    wire N__33122;
    wire N__33119;
    wire N__33114;
    wire N__33107;
    wire N__33104;
    wire N__33099;
    wire N__33094;
    wire N__33091;
    wire N__33090;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33060;
    wire N__33059;
    wire N__33058;
    wire N__33055;
    wire N__33050;
    wire N__33049;
    wire N__33048;
    wire N__33047;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33043;
    wire N__33042;
    wire N__33041;
    wire N__33038;
    wire N__33033;
    wire N__33030;
    wire N__33025;
    wire N__33018;
    wire N__33013;
    wire N__33008;
    wire N__32999;
    wire N__32988;
    wire N__32969;
    wire N__32968;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32936;
    wire N__32935;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32909;
    wire N__32906;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32875;
    wire N__32872;
    wire N__32871;
    wire N__32870;
    wire N__32867;
    wire N__32866;
    wire N__32863;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32831;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32816;
    wire N__32811;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32795;
    wire N__32794;
    wire N__32791;
    wire N__32790;
    wire N__32789;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32759;
    wire N__32756;
    wire N__32749;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32725;
    wire N__32724;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32713;
    wire N__32710;
    wire N__32705;
    wire N__32702;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32670;
    wire N__32667;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32639;
    wire N__32636;
    wire N__32631;
    wire N__32628;
    wire N__32621;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32569;
    wire N__32566;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32435;
    wire N__32432;
    wire N__32431;
    wire N__32430;
    wire N__32427;
    wire N__32426;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32390;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32365;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32357;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32101;
    wire N__32098;
    wire N__32095;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32051;
    wire N__32048;
    wire N__32045;
    wire N__32044;
    wire N__32041;
    wire N__32038;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31916;
    wire N__31913;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31877;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31855;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31847;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31814;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31796;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31785;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31745;
    wire N__31744;
    wire N__31741;
    wire N__31740;
    wire N__31739;
    wire N__31736;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31697;
    wire N__31692;
    wire N__31685;
    wire N__31684;
    wire N__31683;
    wire N__31682;
    wire N__31679;
    wire N__31678;
    wire N__31675;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31647;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31616;
    wire N__31615;
    wire N__31612;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31601;
    wire N__31600;
    wire N__31597;
    wire N__31592;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31546;
    wire N__31543;
    wire N__31540;
    wire N__31539;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31523;
    wire N__31522;
    wire N__31521;
    wire N__31520;
    wire N__31519;
    wire N__31518;
    wire N__31517;
    wire N__31516;
    wire N__31515;
    wire N__31514;
    wire N__31513;
    wire N__31512;
    wire N__31511;
    wire N__31510;
    wire N__31509;
    wire N__31508;
    wire N__31507;
    wire N__31506;
    wire N__31505;
    wire N__31504;
    wire N__31503;
    wire N__31502;
    wire N__31501;
    wire N__31500;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31494;
    wire N__31489;
    wire N__31482;
    wire N__31479;
    wire N__31470;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31448;
    wire N__31433;
    wire N__31432;
    wire N__31431;
    wire N__31430;
    wire N__31429;
    wire N__31428;
    wire N__31427;
    wire N__31426;
    wire N__31425;
    wire N__31424;
    wire N__31423;
    wire N__31422;
    wire N__31421;
    wire N__31418;
    wire N__31415;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31399;
    wire N__31398;
    wire N__31397;
    wire N__31396;
    wire N__31395;
    wire N__31394;
    wire N__31393;
    wire N__31392;
    wire N__31391;
    wire N__31384;
    wire N__31375;
    wire N__31372;
    wire N__31357;
    wire N__31352;
    wire N__31349;
    wire N__31344;
    wire N__31329;
    wire N__31320;
    wire N__31315;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31250;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31235;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31190;
    wire N__31189;
    wire N__31186;
    wire N__31185;
    wire N__31182;
    wire N__31181;
    wire N__31178;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31154;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31118;
    wire N__31117;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31094;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31086;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31063;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31048;
    wire N__31043;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30937;
    wire N__30936;
    wire N__30935;
    wire N__30934;
    wire N__30933;
    wire N__30928;
    wire N__30927;
    wire N__30924;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30872;
    wire N__30871;
    wire N__30870;
    wire N__30869;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30766;
    wire N__30765;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30748;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30703;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30679;
    wire N__30678;
    wire N__30677;
    wire N__30674;
    wire N__30669;
    wire N__30666;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30565;
    wire N__30564;
    wire N__30563;
    wire N__30560;
    wire N__30555;
    wire N__30552;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30505;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30488;
    wire N__30487;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30463;
    wire N__30460;
    wire N__30455;
    wire N__30452;
    wire N__30451;
    wire N__30448;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30434;
    wire N__30431;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30391;
    wire N__30388;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30362;
    wire N__30361;
    wire N__30358;
    wire N__30357;
    wire N__30354;
    wire N__30353;
    wire N__30350;
    wire N__30349;
    wire N__30346;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30324;
    wire N__30319;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30286;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30231;
    wire N__30230;
    wire N__30229;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30043;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30028;
    wire N__30025;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30006;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29971;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29864;
    wire N__29861;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29818;
    wire N__29815;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29744;
    wire N__29741;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29716;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29650;
    wire N__29647;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29630;
    wire N__29629;
    wire N__29626;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29609;
    wire N__29608;
    wire N__29605;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29569;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29518;
    wire N__29517;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29503;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29413;
    wire N__29412;
    wire N__29411;
    wire N__29410;
    wire N__29409;
    wire N__29406;
    wire N__29395;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29363;
    wire N__29360;
    wire N__29355;
    wire N__29352;
    wire N__29345;
    wire N__29344;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29309;
    wire N__29306;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29245;
    wire N__29240;
    wire N__29237;
    wire N__29236;
    wire N__29231;
    wire N__29228;
    wire N__29227;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29207;
    wire N__29204;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29174;
    wire N__29171;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29156;
    wire N__29153;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29141;
    wire N__29138;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29123;
    wire N__29120;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29053;
    wire N__29052;
    wire N__29049;
    wire N__29044;
    wire N__29039;
    wire N__29036;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29018;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28978;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28949;
    wire N__28948;
    wire N__28945;
    wire N__28944;
    wire N__28941;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28923;
    wire N__28918;
    wire N__28915;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28900;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28885;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28843;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28802;
    wire N__28793;
    wire N__28790;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28763;
    wire N__28760;
    wire N__28759;
    wire N__28758;
    wire N__28757;
    wire N__28754;
    wire N__28747;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28729;
    wire N__28726;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28697;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28681;
    wire N__28678;
    wire N__28677;
    wire N__28674;
    wire N__28667;
    wire N__28664;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28660;
    wire N__28659;
    wire N__28658;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28650;
    wire N__28647;
    wire N__28646;
    wire N__28643;
    wire N__28642;
    wire N__28639;
    wire N__28638;
    wire N__28635;
    wire N__28634;
    wire N__28633;
    wire N__28624;
    wire N__28607;
    wire N__28606;
    wire N__28603;
    wire N__28602;
    wire N__28599;
    wire N__28594;
    wire N__28585;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28547;
    wire N__28546;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28523;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28515;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28499;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28477;
    wire N__28472;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28464;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28431;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28396;
    wire N__28393;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28375;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28327;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28303;
    wire N__28302;
    wire N__28301;
    wire N__28300;
    wire N__28299;
    wire N__28298;
    wire N__28297;
    wire N__28296;
    wire N__28295;
    wire N__28294;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28285;
    wire N__28284;
    wire N__28283;
    wire N__28282;
    wire N__28281;
    wire N__28280;
    wire N__28279;
    wire N__28274;
    wire N__28269;
    wire N__28266;
    wire N__28255;
    wire N__28254;
    wire N__28253;
    wire N__28252;
    wire N__28251;
    wire N__28250;
    wire N__28249;
    wire N__28248;
    wire N__28247;
    wire N__28246;
    wire N__28243;
    wire N__28242;
    wire N__28241;
    wire N__28230;
    wire N__28221;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28205;
    wire N__28196;
    wire N__28183;
    wire N__28178;
    wire N__28173;
    wire N__28170;
    wire N__28157;
    wire N__28156;
    wire N__28155;
    wire N__28154;
    wire N__28153;
    wire N__28152;
    wire N__28151;
    wire N__28150;
    wire N__28149;
    wire N__28148;
    wire N__28147;
    wire N__28146;
    wire N__28145;
    wire N__28144;
    wire N__28133;
    wire N__28132;
    wire N__28131;
    wire N__28130;
    wire N__28129;
    wire N__28128;
    wire N__28127;
    wire N__28126;
    wire N__28125;
    wire N__28124;
    wire N__28123;
    wire N__28122;
    wire N__28121;
    wire N__28108;
    wire N__28103;
    wire N__28102;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28084;
    wire N__28083;
    wire N__28074;
    wire N__28063;
    wire N__28058;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28032;
    wire N__28025;
    wire N__28018;
    wire N__28007;
    wire N__28006;
    wire N__28005;
    wire N__28004;
    wire N__28003;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27987;
    wire N__27986;
    wire N__27985;
    wire N__27982;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27971;
    wire N__27970;
    wire N__27969;
    wire N__27968;
    wire N__27967;
    wire N__27966;
    wire N__27965;
    wire N__27964;
    wire N__27959;
    wire N__27948;
    wire N__27939;
    wire N__27928;
    wire N__27923;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27915;
    wire N__27914;
    wire N__27907;
    wire N__27904;
    wire N__27903;
    wire N__27900;
    wire N__27895;
    wire N__27890;
    wire N__27887;
    wire N__27886;
    wire N__27885;
    wire N__27884;
    wire N__27883;
    wire N__27882;
    wire N__27881;
    wire N__27880;
    wire N__27879;
    wire N__27874;
    wire N__27871;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27820;
    wire N__27813;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27793;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27748;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27716;
    wire N__27713;
    wire N__27708;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27650;
    wire N__27649;
    wire N__27646;
    wire N__27645;
    wire N__27642;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27575;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27457;
    wire N__27454;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27443;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27428;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27406;
    wire N__27403;
    wire N__27402;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27301;
    wire N__27298;
    wire N__27297;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27276;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27219;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27208;
    wire N__27205;
    wire N__27200;
    wire N__27197;
    wire N__27192;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26938;
    wire N__26937;
    wire N__26936;
    wire N__26935;
    wire N__26934;
    wire N__26933;
    wire N__26932;
    wire N__26931;
    wire N__26930;
    wire N__26929;
    wire N__26928;
    wire N__26927;
    wire N__26926;
    wire N__26925;
    wire N__26924;
    wire N__26923;
    wire N__26922;
    wire N__26921;
    wire N__26920;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26916;
    wire N__26915;
    wire N__26914;
    wire N__26913;
    wire N__26912;
    wire N__26911;
    wire N__26910;
    wire N__26901;
    wire N__26892;
    wire N__26883;
    wire N__26874;
    wire N__26869;
    wire N__26860;
    wire N__26851;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26806;
    wire N__26803;
    wire N__26798;
    wire N__26795;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26765;
    wire N__26764;
    wire N__26763;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26751;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26669;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26634;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26611;
    wire N__26608;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26593;
    wire N__26588;
    wire N__26585;
    wire N__26584;
    wire N__26579;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26557;
    wire N__26554;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26524;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26487;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26471;
    wire N__26468;
    wire N__26467;
    wire N__26466;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26450;
    wire N__26447;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26432;
    wire N__26429;
    wire N__26428;
    wire N__26427;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26411;
    wire N__26408;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26400;
    wire N__26395;
    wire N__26392;
    wire N__26389;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26377;
    wire N__26374;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26359;
    wire N__26354;
    wire N__26351;
    wire N__26350;
    wire N__26345;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26330;
    wire N__26327;
    wire N__26326;
    wire N__26323;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26290;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26274;
    wire N__26267;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26256;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26240;
    wire N__26237;
    wire N__26236;
    wire N__26235;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26214;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26198;
    wire N__26195;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26183;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26168;
    wire N__26165;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26157;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26137;
    wire N__26136;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26120;
    wire N__26117;
    wire N__26116;
    wire N__26111;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26089;
    wire N__26086;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26056;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26033;
    wire N__26030;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26006;
    wire N__26003;
    wire N__26002;
    wire N__26001;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25978;
    wire N__25975;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25960;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25939;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25925;
    wire N__25922;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25859;
    wire N__25856;
    wire N__25855;
    wire N__25854;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25017;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24989;
    wire N__24980;
    wire N__24977;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24969;
    wire N__24966;
    wire N__24965;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24944;
    wire N__24935;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24926;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24900;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24886;
    wire N__24885;
    wire N__24884;
    wire N__24881;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24860;
    wire N__24857;
    wire N__24848;
    wire N__24845;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24833;
    wire N__24832;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24815;
    wire N__24814;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24761;
    wire N__24756;
    wire N__24751;
    wire N__24746;
    wire N__24745;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24728;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24688;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24598;
    wire N__24597;
    wire N__24596;
    wire N__24595;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24571;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24559;
    wire N__24554;
    wire N__24551;
    wire N__24550;
    wire N__24547;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24520;
    wire N__24517;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24502;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24473;
    wire N__24472;
    wire N__24471;
    wire N__24468;
    wire N__24463;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24431;
    wire N__24428;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24416;
    wire N__24415;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24391;
    wire N__24386;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24361;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24337;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24304;
    wire N__24303;
    wire N__24300;
    wire N__24295;
    wire N__24290;
    wire N__24287;
    wire N__24286;
    wire N__24285;
    wire N__24284;
    wire N__24281;
    wire N__24276;
    wire N__24273;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24241;
    wire N__24240;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24224;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23872;
    wire N__23869;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23852;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23743;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23704;
    wire N__23703;
    wire N__23702;
    wire N__23699;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23667;
    wire N__23660;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23648;
    wire N__23645;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23630;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23579;
    wire N__23576;
    wire N__23575;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23543;
    wire N__23542;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23516;
    wire N__23515;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23496;
    wire N__23493;
    wire N__23488;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22831;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22801;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22724;
    wire N__22721;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22673;
    wire N__22670;
    wire N__22669;
    wire N__22668;
    wire N__22667;
    wire N__22662;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22641;
    wire N__22638;
    wire N__22633;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22601;
    wire N__22598;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22573;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22558;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22495;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22477;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22429;
    wire N__22428;
    wire N__22425;
    wire N__22420;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22392;
    wire N__22389;
    wire N__22384;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22340;
    wire N__22337;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22255;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22240;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22209;
    wire N__22208;
    wire N__22205;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22177;
    wire N__22176;
    wire N__22173;
    wire N__22168;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22156;
    wire N__22155;
    wire N__22152;
    wire N__22147;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22132;
    wire N__22131;
    wire N__22128;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22039;
    wire N__22038;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22031;
    wire N__22024;
    wire N__22019;
    wire N__22016;
    wire N__22011;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21922;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21877;
    wire N__21874;
    wire N__21873;
    wire N__21872;
    wire N__21871;
    wire N__21870;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21864;
    wire N__21859;
    wire N__21854;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21836;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21748;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21673;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21411;
    wire N__21410;
    wire N__21409;
    wire N__21408;
    wire N__21407;
    wire N__21406;
    wire N__21405;
    wire N__21404;
    wire N__21399;
    wire N__21396;
    wire N__21391;
    wire N__21388;
    wire N__21379;
    wire N__21372;
    wire N__21369;
    wire N__21364;
    wire N__21359;
    wire N__21358;
    wire N__21357;
    wire N__21356;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21343;
    wire N__21334;
    wire N__21331;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21323;
    wire N__21318;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21298;
    wire N__21295;
    wire N__21290;
    wire N__21289;
    wire N__21288;
    wire N__21287;
    wire N__21286;
    wire N__21283;
    wire N__21274;
    wire N__21273;
    wire N__21270;
    wire N__21269;
    wire N__21266;
    wire N__21265;
    wire N__21264;
    wire N__21263;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21254;
    wire N__21253;
    wire N__21252;
    wire N__21251;
    wire N__21250;
    wire N__21249;
    wire N__21248;
    wire N__21247;
    wire N__21246;
    wire N__21245;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21233;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21213;
    wire N__21196;
    wire N__21193;
    wire N__21186;
    wire N__21179;
    wire N__21178;
    wire N__21177;
    wire N__21176;
    wire N__21175;
    wire N__21174;
    wire N__21173;
    wire N__21172;
    wire N__21171;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21137;
    wire N__21134;
    wire N__21129;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21094;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21070;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21037;
    wire N__21034;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21010;
    wire N__21007;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20916;
    wire N__20915;
    wire N__20914;
    wire N__20913;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20894;
    wire N__20889;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20855;
    wire N__20854;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20750;
    wire N__20749;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20714;
    wire N__20713;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20693;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20675;
    wire N__20672;
    wire N__20671;
    wire N__20668;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20651;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20639;
    wire N__20638;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20617;
    wire N__20616;
    wire N__20613;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20601;
    wire N__20600;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20582;
    wire N__20579;
    wire N__20568;
    wire N__20565;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20338;
    wire N__20337;
    wire N__20334;
    wire N__20329;
    wire N__20324;
    wire N__20323;
    wire N__20320;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20302;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20266;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20249;
    wire N__20248;
    wire N__20247;
    wire N__20244;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20215;
    wire N__20210;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20075;
    wire N__20066;
    wire N__20063;
    wire N__20062;
    wire N__20059;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20042;
    wire N__20039;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20027;
    wire N__20024;
    wire N__20023;
    wire N__20022;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19991;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19976;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19961;
    wire N__19960;
    wire N__19959;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19825;
    wire N__19822;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19807;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19786;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19558;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19353;
    wire N__19350;
    wire N__19349;
    wire N__19346;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19326;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire bfn_1_13_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_1_17_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_1_18_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_1_19_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire N_34_i_i;
    wire rgb_drv_RNOZ0;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.N_168_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_166 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_166_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_162 ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.N_167 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_6;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ;
    wire pwm_duty_input_8;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire bfn_2_13_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire bfn_2_14_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire bfn_2_16_0_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire bfn_2_17_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_3_10_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.N_17 ;
    wire N_19_1;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_4_9_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_4_10_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire il_max_comp2_c;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire il_max_comp2_D1;
    wire il_min_comp2_c;
    wire il_min_comp2_D1;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire bfn_7_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire bfn_7_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire bfn_7_13_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire bfn_7_14_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire bfn_7_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_7_16_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_7_17_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire \delay_measurement_inst.N_34 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_ ;
    wire \delay_measurement_inst.N_32 ;
    wire \delay_measurement_inst.N_35 ;
    wire \delay_measurement_inst.N_43 ;
    wire il_max_comp1_c;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_74_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.N_71 ;
    wire \current_shift_inst.PI_CTRL.N_75_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire s4_phy_c;
    wire \delay_measurement_inst.N_31 ;
    wire \delay_measurement_inst.N_40 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt14_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_4_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0 ;
    wire \delay_measurement_inst.un1_elapsed_time_hc_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ;
    wire \delay_measurement_inst.N_30_cascade_ ;
    wire \delay_measurement_inst.N_37 ;
    wire \delay_measurement_inst.delay_hc_timer.N_302_i ;
    wire \delay_measurement_inst.N_36 ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire il_min_comp2_D2;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_72 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_9_14_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire bfn_9_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_9_16_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt30_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt14_0 ;
    wire \delay_measurement_inst.N_41 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire bfn_9_19_0_;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_9_20_0_;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire bfn_9_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_9_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_302_i_g ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.N_52 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire il_min_comp1_c;
    wire il_max_comp1_D1;
    wire il_min_comp1_D1;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_16 ;
    wire bfn_10_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire bfn_10_11_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_10_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire bfn_10_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_10_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_10_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_10_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_10_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_10_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.N_39_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_27 ;
    wire s3_phy_c;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_11_8_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire bfn_11_9_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire bfn_11_10_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire bfn_11_11_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.N_74 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.N_33_cascade_ ;
    wire \delay_measurement_inst.N_38 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.N_303_i ;
    wire \delay_measurement_inst.N_28 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire measured_delay_hc_25;
    wire measured_delay_hc_24;
    wire measured_delay_hc_26;
    wire measured_delay_hc_23;
    wire measured_delay_hc_28;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.N_51 ;
    wire measured_delay_hc_27;
    wire \delay_measurement_inst.N_25 ;
    wire \delay_measurement_inst.delay_tr_timer.N_304_i ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire delay_tr_d2;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.N_59 ;
    wire \delay_measurement_inst.N_270 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_12_10_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire bfn_12_11_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire bfn_12_13_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_12_14_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_12_15_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire measured_delay_hc_14;
    wire \phase_controller_inst1.stoper_hc.un1_startlt8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire measured_delay_hc_19;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire measured_delay_hc_17;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3 ;
    wire measured_delay_hc_20;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.N_29_cascade_ ;
    wire measured_delay_hc_6;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6 ;
    wire measured_delay_hc_21;
    wire \delay_measurement_inst.N_42 ;
    wire measured_delay_hc_18;
    wire \delay_measurement_inst.N_26 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \delay_measurement_inst.N_27 ;
    wire \delay_measurement_inst.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.N_53 ;
    wire measured_delay_hc_29;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3 ;
    wire \delay_measurement_inst.N_54 ;
    wire measured_delay_hc_30;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire delay_hc_d2;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7 ;
    wire \delay_measurement_inst.N_299 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire bfn_13_12_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire bfn_13_13_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_16 ;
    wire bfn_13_14_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire measured_delay_hc_4;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire measured_delay_hc_5;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire measured_delay_hc_16;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire measured_delay_hc_1;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_start ;
    wire measured_delay_hc_3;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire measured_delay_hc_7;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire measured_delay_hc_8;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ;
    wire measured_delay_hc_0;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ;
    wire measured_delay_hc_13;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire measured_delay_hc_15;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt30 ;
    wire measured_delay_hc_2;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire il_max_comp1_D2;
    wire state_ns_i_a3_1;
    wire measured_delay_hc_12;
    wire measured_delay_hc_11;
    wire measured_delay_hc_9;
    wire measured_delay_hc_10;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire \delay_measurement_inst.delay_hc_reg3lt31_0 ;
    wire measured_delay_hc_22;
    wire state_3;
    wire s1_phy_c;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_181_i ;
    wire s2_phy_c;
    wire \phase_controller_inst2.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_14_6_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_14_7_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_17 ;
    wire bfn_14_8_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire measured_delay_tr_5;
    wire measured_delay_tr_3;
    wire \phase_controller_inst1.stoper_tr.N_248 ;
    wire measured_delay_tr_1;
    wire measured_delay_tr_11;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ;
    wire measured_delay_tr_6;
    wire measured_delay_tr_2;
    wire \phase_controller_inst1.stoper_tr.N_55 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire red_c_i;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hc_RNO_0_0_cascade_ ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire il_max_comp2_D2;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire measured_delay_hc_31;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.time_passed11 ;
    wire \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire bfn_15_2_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire bfn_15_3_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire bfn_15_4_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.N_290 ;
    wire \delay_measurement_inst.N_325 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire measured_delay_tr_10;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ;
    wire measured_delay_tr_4;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.time_passed11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ;
    wire measured_delay_tr_19;
    wire measured_delay_tr_12;
    wire measured_delay_tr_14;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ;
    wire measured_delay_tr_13;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ;
    wire measured_delay_tr_15;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_10_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_11_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_15_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire measured_delay_tr_17;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire measured_delay_tr_18;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire measured_delay_tr_7;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i ;
    wire \delay_measurement_inst.N_267 ;
    wire measured_delay_tr_8;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.N_1318_i ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire bfn_15_18_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_15_19_0_;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_15_20_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_15_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_15_23_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_15_24_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire bfn_15_25_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_15_26_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_15_27_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_15_28_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_181_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ;
    wire \delay_measurement_inst.N_265 ;
    wire \delay_measurement_inst.delay_tr_timer.N_287_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_16_7_0_;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_reg3lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_reg3lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_16_8_0_;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_reg3lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_reg3lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_16_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_16_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_16_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire bfn_16_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_16_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire bfn_16_14_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un4_control_input_0_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire measured_delay_tr_16;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire bfn_17_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_17_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_17_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_305_i ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_17_19_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.N_304_i_g ;
    wire start_stop_c;
    wire phase_controller_inst1_state_4;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire bfn_18_13_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_18_14_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_18_15_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_18_16_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \current_shift_inst.timer_s1.N_180_i_g ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__24662),
            .RESETB(N__35913),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__46031),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__46024),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__21250,N__21176,N__21248,N__21175,N__21249,N__21174,N__21251,N__21171,N__21244,N__21170,N__21245,N__21172,N__21246,N__21173,N__21247}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__46030,N__46027,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__46025,N__46029,N__46026,N__46028}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__45857),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__45890),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__21261,N__21264,N__21262,N__21265,N__21263,N__20319,N__20265,N__21033,N__20295,N__21006,N__20209,N__20249,N__19976,N__19991,N__20006}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__45896,N__45893,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__45891,N__45895,N__45892,N__45894}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__49947),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__49949),
            .DIN(N__49948),
            .DOUT(N__49947),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__49949),
            .PADOUT(N__49948),
            .PADIN(N__49947),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__49938),
            .DIN(N__49937),
            .DOUT(N__49936),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__49938),
            .PADOUT(N__49937),
            .PADIN(N__49936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__49929),
            .DIN(N__49928),
            .DOUT(N__49927),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__49929),
            .PADOUT(N__49928),
            .PADIN(N__49927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__49920),
            .DIN(N__49919),
            .DOUT(N__49918),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__49920),
            .PADOUT(N__49919),
            .PADIN(N__49918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21893),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__49911),
            .DIN(N__49910),
            .DOUT(N__49909),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__49911),
            .PADOUT(N__49910),
            .PADIN(N__49909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__49902),
            .DIN(N__49901),
            .DOUT(N__49900),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__49902),
            .PADOUT(N__49901),
            .PADIN(N__49900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__49893),
            .DIN(N__49892),
            .DOUT(N__49891),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__49893),
            .PADOUT(N__49892),
            .PADIN(N__49891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__49884),
            .DIN(N__49883),
            .DOUT(N__49882),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__49884),
            .PADOUT(N__49883),
            .PADIN(N__49882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__49875),
            .DIN(N__49874),
            .DOUT(N__49873),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__49875),
            .PADOUT(N__49874),
            .PADIN(N__49873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__49866),
            .DIN(N__49865),
            .DOUT(N__49864),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__49866),
            .PADOUT(N__49865),
            .PADIN(N__49864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34574),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__49857),
            .DIN(N__49856),
            .DOUT(N__49855),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__49857),
            .PADOUT(N__49856),
            .PADIN(N__49855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23249),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__49848),
            .DIN(N__49847),
            .DOUT(N__49846),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__49848),
            .PADOUT(N__49847),
            .PADIN(N__49846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__49839),
            .DIN(N__49838),
            .DOUT(N__49837),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__49839),
            .PADOUT(N__49838),
            .PADIN(N__49837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11854 (
            .O(N__49820),
            .I(N__49817));
    LocalMux I__11853 (
            .O(N__49817),
            .I(N__49814));
    Odrv12 I__11852 (
            .O(N__49814),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__11851 (
            .O(N__49811),
            .I(N__49808));
    LocalMux I__11850 (
            .O(N__49808),
            .I(N__49805));
    Odrv12 I__11849 (
            .O(N__49805),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__11848 (
            .O(N__49802),
            .I(N__49799));
    LocalMux I__11847 (
            .O(N__49799),
            .I(N__49796));
    Span4Mux_h I__11846 (
            .O(N__49796),
            .I(N__49793));
    Odrv4 I__11845 (
            .O(N__49793),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__11844 (
            .O(N__49790),
            .I(N__49787));
    LocalMux I__11843 (
            .O(N__49787),
            .I(N__49772));
    InMux I__11842 (
            .O(N__49786),
            .I(N__49767));
    InMux I__11841 (
            .O(N__49785),
            .I(N__49767));
    InMux I__11840 (
            .O(N__49784),
            .I(N__49758));
    InMux I__11839 (
            .O(N__49783),
            .I(N__49729));
    InMux I__11838 (
            .O(N__49782),
            .I(N__49716));
    InMux I__11837 (
            .O(N__49781),
            .I(N__49716));
    InMux I__11836 (
            .O(N__49780),
            .I(N__49716));
    InMux I__11835 (
            .O(N__49779),
            .I(N__49716));
    InMux I__11834 (
            .O(N__49778),
            .I(N__49716));
    InMux I__11833 (
            .O(N__49777),
            .I(N__49716));
    InMux I__11832 (
            .O(N__49776),
            .I(N__49711));
    InMux I__11831 (
            .O(N__49775),
            .I(N__49711));
    Span4Mux_v I__11830 (
            .O(N__49772),
            .I(N__49702));
    LocalMux I__11829 (
            .O(N__49767),
            .I(N__49702));
    InMux I__11828 (
            .O(N__49766),
            .I(N__49699));
    InMux I__11827 (
            .O(N__49765),
            .I(N__49688));
    InMux I__11826 (
            .O(N__49764),
            .I(N__49688));
    InMux I__11825 (
            .O(N__49763),
            .I(N__49688));
    InMux I__11824 (
            .O(N__49762),
            .I(N__49688));
    InMux I__11823 (
            .O(N__49761),
            .I(N__49688));
    LocalMux I__11822 (
            .O(N__49758),
            .I(N__49685));
    InMux I__11821 (
            .O(N__49757),
            .I(N__49670));
    InMux I__11820 (
            .O(N__49756),
            .I(N__49670));
    InMux I__11819 (
            .O(N__49755),
            .I(N__49670));
    InMux I__11818 (
            .O(N__49754),
            .I(N__49670));
    InMux I__11817 (
            .O(N__49753),
            .I(N__49670));
    InMux I__11816 (
            .O(N__49752),
            .I(N__49670));
    InMux I__11815 (
            .O(N__49751),
            .I(N__49670));
    InMux I__11814 (
            .O(N__49750),
            .I(N__49665));
    InMux I__11813 (
            .O(N__49749),
            .I(N__49665));
    InMux I__11812 (
            .O(N__49748),
            .I(N__49660));
    InMux I__11811 (
            .O(N__49747),
            .I(N__49660));
    InMux I__11810 (
            .O(N__49746),
            .I(N__49655));
    InMux I__11809 (
            .O(N__49745),
            .I(N__49655));
    InMux I__11808 (
            .O(N__49744),
            .I(N__49646));
    InMux I__11807 (
            .O(N__49743),
            .I(N__49646));
    InMux I__11806 (
            .O(N__49742),
            .I(N__49646));
    InMux I__11805 (
            .O(N__49741),
            .I(N__49646));
    InMux I__11804 (
            .O(N__49740),
            .I(N__49636));
    InMux I__11803 (
            .O(N__49739),
            .I(N__49636));
    InMux I__11802 (
            .O(N__49738),
            .I(N__49636));
    InMux I__11801 (
            .O(N__49737),
            .I(N__49636));
    InMux I__11800 (
            .O(N__49736),
            .I(N__49625));
    InMux I__11799 (
            .O(N__49735),
            .I(N__49625));
    InMux I__11798 (
            .O(N__49734),
            .I(N__49625));
    InMux I__11797 (
            .O(N__49733),
            .I(N__49625));
    InMux I__11796 (
            .O(N__49732),
            .I(N__49625));
    LocalMux I__11795 (
            .O(N__49729),
            .I(N__49610));
    LocalMux I__11794 (
            .O(N__49716),
            .I(N__49610));
    LocalMux I__11793 (
            .O(N__49711),
            .I(N__49610));
    InMux I__11792 (
            .O(N__49710),
            .I(N__49607));
    InMux I__11791 (
            .O(N__49709),
            .I(N__49604));
    InMux I__11790 (
            .O(N__49708),
            .I(N__49599));
    InMux I__11789 (
            .O(N__49707),
            .I(N__49599));
    Span4Mux_v I__11788 (
            .O(N__49702),
            .I(N__49596));
    LocalMux I__11787 (
            .O(N__49699),
            .I(N__49591));
    LocalMux I__11786 (
            .O(N__49688),
            .I(N__49591));
    Span4Mux_v I__11785 (
            .O(N__49685),
            .I(N__49582));
    LocalMux I__11784 (
            .O(N__49670),
            .I(N__49582));
    LocalMux I__11783 (
            .O(N__49665),
            .I(N__49570));
    LocalMux I__11782 (
            .O(N__49660),
            .I(N__49570));
    LocalMux I__11781 (
            .O(N__49655),
            .I(N__49570));
    LocalMux I__11780 (
            .O(N__49646),
            .I(N__49567));
    CascadeMux I__11779 (
            .O(N__49645),
            .I(N__49562));
    LocalMux I__11778 (
            .O(N__49636),
            .I(N__49556));
    LocalMux I__11777 (
            .O(N__49625),
            .I(N__49556));
    InMux I__11776 (
            .O(N__49624),
            .I(N__49539));
    InMux I__11775 (
            .O(N__49623),
            .I(N__49539));
    InMux I__11774 (
            .O(N__49622),
            .I(N__49539));
    InMux I__11773 (
            .O(N__49621),
            .I(N__49539));
    InMux I__11772 (
            .O(N__49620),
            .I(N__49539));
    InMux I__11771 (
            .O(N__49619),
            .I(N__49539));
    InMux I__11770 (
            .O(N__49618),
            .I(N__49539));
    InMux I__11769 (
            .O(N__49617),
            .I(N__49539));
    Span4Mux_v I__11768 (
            .O(N__49610),
            .I(N__49534));
    LocalMux I__11767 (
            .O(N__49607),
            .I(N__49534));
    LocalMux I__11766 (
            .O(N__49604),
            .I(N__49529));
    LocalMux I__11765 (
            .O(N__49599),
            .I(N__49529));
    Span4Mux_h I__11764 (
            .O(N__49596),
            .I(N__49526));
    Span12Mux_s11_h I__11763 (
            .O(N__49591),
            .I(N__49523));
    InMux I__11762 (
            .O(N__49590),
            .I(N__49514));
    InMux I__11761 (
            .O(N__49589),
            .I(N__49514));
    InMux I__11760 (
            .O(N__49588),
            .I(N__49514));
    InMux I__11759 (
            .O(N__49587),
            .I(N__49514));
    Span4Mux_h I__11758 (
            .O(N__49582),
            .I(N__49511));
    InMux I__11757 (
            .O(N__49581),
            .I(N__49508));
    InMux I__11756 (
            .O(N__49580),
            .I(N__49499));
    InMux I__11755 (
            .O(N__49579),
            .I(N__49499));
    InMux I__11754 (
            .O(N__49578),
            .I(N__49499));
    InMux I__11753 (
            .O(N__49577),
            .I(N__49499));
    Span4Mux_h I__11752 (
            .O(N__49570),
            .I(N__49494));
    Span4Mux_h I__11751 (
            .O(N__49567),
            .I(N__49494));
    InMux I__11750 (
            .O(N__49566),
            .I(N__49485));
    InMux I__11749 (
            .O(N__49565),
            .I(N__49485));
    InMux I__11748 (
            .O(N__49562),
            .I(N__49485));
    InMux I__11747 (
            .O(N__49561),
            .I(N__49485));
    Span4Mux_v I__11746 (
            .O(N__49556),
            .I(N__49476));
    LocalMux I__11745 (
            .O(N__49539),
            .I(N__49476));
    Span4Mux_h I__11744 (
            .O(N__49534),
            .I(N__49476));
    Span4Mux_v I__11743 (
            .O(N__49529),
            .I(N__49476));
    Odrv4 I__11742 (
            .O(N__49526),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__11741 (
            .O(N__49523),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11740 (
            .O(N__49514),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11739 (
            .O(N__49511),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11738 (
            .O(N__49508),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11737 (
            .O(N__49499),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11736 (
            .O(N__49494),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11735 (
            .O(N__49485),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11734 (
            .O(N__49476),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__11733 (
            .O(N__49457),
            .I(N__49451));
    CascadeMux I__11732 (
            .O(N__49456),
            .I(N__49447));
    CascadeMux I__11731 (
            .O(N__49455),
            .I(N__49444));
    CascadeMux I__11730 (
            .O(N__49454),
            .I(N__49440));
    InMux I__11729 (
            .O(N__49451),
            .I(N__49436));
    CascadeMux I__11728 (
            .O(N__49450),
            .I(N__49424));
    InMux I__11727 (
            .O(N__49447),
            .I(N__49420));
    InMux I__11726 (
            .O(N__49444),
            .I(N__49417));
    InMux I__11725 (
            .O(N__49443),
            .I(N__49414));
    InMux I__11724 (
            .O(N__49440),
            .I(N__49409));
    InMux I__11723 (
            .O(N__49439),
            .I(N__49409));
    LocalMux I__11722 (
            .O(N__49436),
            .I(N__49406));
    CascadeMux I__11721 (
            .O(N__49435),
            .I(N__49403));
    CascadeMux I__11720 (
            .O(N__49434),
            .I(N__49397));
    CascadeMux I__11719 (
            .O(N__49433),
            .I(N__49385));
    CascadeMux I__11718 (
            .O(N__49432),
            .I(N__49382));
    CascadeMux I__11717 (
            .O(N__49431),
            .I(N__49374));
    CascadeMux I__11716 (
            .O(N__49430),
            .I(N__49371));
    CascadeMux I__11715 (
            .O(N__49429),
            .I(N__49366));
    CascadeMux I__11714 (
            .O(N__49428),
            .I(N__49363));
    InMux I__11713 (
            .O(N__49427),
            .I(N__49342));
    InMux I__11712 (
            .O(N__49424),
            .I(N__49342));
    InMux I__11711 (
            .O(N__49423),
            .I(N__49342));
    LocalMux I__11710 (
            .O(N__49420),
            .I(N__49337));
    LocalMux I__11709 (
            .O(N__49417),
            .I(N__49337));
    LocalMux I__11708 (
            .O(N__49414),
            .I(N__49332));
    LocalMux I__11707 (
            .O(N__49409),
            .I(N__49332));
    Span4Mux_h I__11706 (
            .O(N__49406),
            .I(N__49329));
    InMux I__11705 (
            .O(N__49403),
            .I(N__49318));
    InMux I__11704 (
            .O(N__49402),
            .I(N__49318));
    InMux I__11703 (
            .O(N__49401),
            .I(N__49318));
    InMux I__11702 (
            .O(N__49400),
            .I(N__49318));
    InMux I__11701 (
            .O(N__49397),
            .I(N__49318));
    CascadeMux I__11700 (
            .O(N__49396),
            .I(N__49315));
    CascadeMux I__11699 (
            .O(N__49395),
            .I(N__49312));
    CascadeMux I__11698 (
            .O(N__49394),
            .I(N__49305));
    CascadeMux I__11697 (
            .O(N__49393),
            .I(N__49302));
    CascadeMux I__11696 (
            .O(N__49392),
            .I(N__49299));
    CascadeMux I__11695 (
            .O(N__49391),
            .I(N__49296));
    CascadeMux I__11694 (
            .O(N__49390),
            .I(N__49293));
    CascadeMux I__11693 (
            .O(N__49389),
            .I(N__49289));
    CascadeMux I__11692 (
            .O(N__49388),
            .I(N__49286));
    InMux I__11691 (
            .O(N__49385),
            .I(N__49267));
    InMux I__11690 (
            .O(N__49382),
            .I(N__49267));
    CascadeMux I__11689 (
            .O(N__49381),
            .I(N__49263));
    CascadeMux I__11688 (
            .O(N__49380),
            .I(N__49260));
    CascadeMux I__11687 (
            .O(N__49379),
            .I(N__49257));
    CascadeMux I__11686 (
            .O(N__49378),
            .I(N__49251));
    InMux I__11685 (
            .O(N__49377),
            .I(N__49243));
    InMux I__11684 (
            .O(N__49374),
            .I(N__49243));
    InMux I__11683 (
            .O(N__49371),
            .I(N__49236));
    InMux I__11682 (
            .O(N__49370),
            .I(N__49236));
    InMux I__11681 (
            .O(N__49369),
            .I(N__49236));
    InMux I__11680 (
            .O(N__49366),
            .I(N__49231));
    InMux I__11679 (
            .O(N__49363),
            .I(N__49231));
    CascadeMux I__11678 (
            .O(N__49362),
            .I(N__49228));
    CascadeMux I__11677 (
            .O(N__49361),
            .I(N__49225));
    CascadeMux I__11676 (
            .O(N__49360),
            .I(N__49221));
    CascadeMux I__11675 (
            .O(N__49359),
            .I(N__49217));
    CascadeMux I__11674 (
            .O(N__49358),
            .I(N__49213));
    CascadeMux I__11673 (
            .O(N__49357),
            .I(N__49209));
    CascadeMux I__11672 (
            .O(N__49356),
            .I(N__49205));
    CascadeMux I__11671 (
            .O(N__49355),
            .I(N__49192));
    CascadeMux I__11670 (
            .O(N__49354),
            .I(N__49188));
    CascadeMux I__11669 (
            .O(N__49353),
            .I(N__49184));
    CascadeMux I__11668 (
            .O(N__49352),
            .I(N__49180));
    CascadeMux I__11667 (
            .O(N__49351),
            .I(N__49175));
    CascadeMux I__11666 (
            .O(N__49350),
            .I(N__49171));
    CascadeMux I__11665 (
            .O(N__49349),
            .I(N__49167));
    LocalMux I__11664 (
            .O(N__49342),
            .I(N__49164));
    Span4Mux_v I__11663 (
            .O(N__49337),
            .I(N__49159));
    Span4Mux_v I__11662 (
            .O(N__49332),
            .I(N__49159));
    Span4Mux_h I__11661 (
            .O(N__49329),
            .I(N__49154));
    LocalMux I__11660 (
            .O(N__49318),
            .I(N__49154));
    InMux I__11659 (
            .O(N__49315),
            .I(N__49137));
    InMux I__11658 (
            .O(N__49312),
            .I(N__49137));
    InMux I__11657 (
            .O(N__49311),
            .I(N__49137));
    InMux I__11656 (
            .O(N__49310),
            .I(N__49137));
    InMux I__11655 (
            .O(N__49309),
            .I(N__49137));
    InMux I__11654 (
            .O(N__49308),
            .I(N__49137));
    InMux I__11653 (
            .O(N__49305),
            .I(N__49137));
    InMux I__11652 (
            .O(N__49302),
            .I(N__49137));
    InMux I__11651 (
            .O(N__49299),
            .I(N__49128));
    InMux I__11650 (
            .O(N__49296),
            .I(N__49128));
    InMux I__11649 (
            .O(N__49293),
            .I(N__49128));
    InMux I__11648 (
            .O(N__49292),
            .I(N__49128));
    InMux I__11647 (
            .O(N__49289),
            .I(N__49123));
    InMux I__11646 (
            .O(N__49286),
            .I(N__49123));
    CascadeMux I__11645 (
            .O(N__49285),
            .I(N__49120));
    CascadeMux I__11644 (
            .O(N__49284),
            .I(N__49117));
    CascadeMux I__11643 (
            .O(N__49283),
            .I(N__49114));
    CascadeMux I__11642 (
            .O(N__49282),
            .I(N__49111));
    CascadeMux I__11641 (
            .O(N__49281),
            .I(N__49107));
    CascadeMux I__11640 (
            .O(N__49280),
            .I(N__49100));
    CascadeMux I__11639 (
            .O(N__49279),
            .I(N__49096));
    CascadeMux I__11638 (
            .O(N__49278),
            .I(N__49092));
    CascadeMux I__11637 (
            .O(N__49277),
            .I(N__49088));
    CascadeMux I__11636 (
            .O(N__49276),
            .I(N__49084));
    CascadeMux I__11635 (
            .O(N__49275),
            .I(N__49081));
    CascadeMux I__11634 (
            .O(N__49274),
            .I(N__49077));
    CascadeMux I__11633 (
            .O(N__49273),
            .I(N__49073));
    CascadeMux I__11632 (
            .O(N__49272),
            .I(N__49069));
    LocalMux I__11631 (
            .O(N__49267),
            .I(N__49065));
    InMux I__11630 (
            .O(N__49266),
            .I(N__49060));
    InMux I__11629 (
            .O(N__49263),
            .I(N__49060));
    InMux I__11628 (
            .O(N__49260),
            .I(N__49055));
    InMux I__11627 (
            .O(N__49257),
            .I(N__49055));
    InMux I__11626 (
            .O(N__49256),
            .I(N__49040));
    InMux I__11625 (
            .O(N__49255),
            .I(N__49040));
    InMux I__11624 (
            .O(N__49254),
            .I(N__49040));
    InMux I__11623 (
            .O(N__49251),
            .I(N__49040));
    InMux I__11622 (
            .O(N__49250),
            .I(N__49040));
    InMux I__11621 (
            .O(N__49249),
            .I(N__49040));
    InMux I__11620 (
            .O(N__49248),
            .I(N__49040));
    LocalMux I__11619 (
            .O(N__49243),
            .I(N__49035));
    LocalMux I__11618 (
            .O(N__49236),
            .I(N__49035));
    LocalMux I__11617 (
            .O(N__49231),
            .I(N__49032));
    InMux I__11616 (
            .O(N__49228),
            .I(N__49021));
    InMux I__11615 (
            .O(N__49225),
            .I(N__49021));
    InMux I__11614 (
            .O(N__49224),
            .I(N__49021));
    InMux I__11613 (
            .O(N__49221),
            .I(N__49021));
    InMux I__11612 (
            .O(N__49220),
            .I(N__49021));
    InMux I__11611 (
            .O(N__49217),
            .I(N__49004));
    InMux I__11610 (
            .O(N__49216),
            .I(N__49004));
    InMux I__11609 (
            .O(N__49213),
            .I(N__49004));
    InMux I__11608 (
            .O(N__49212),
            .I(N__49004));
    InMux I__11607 (
            .O(N__49209),
            .I(N__49004));
    InMux I__11606 (
            .O(N__49208),
            .I(N__49004));
    InMux I__11605 (
            .O(N__49205),
            .I(N__49004));
    InMux I__11604 (
            .O(N__49204),
            .I(N__49004));
    CascadeMux I__11603 (
            .O(N__49203),
            .I(N__49001));
    CascadeMux I__11602 (
            .O(N__49202),
            .I(N__48998));
    CascadeMux I__11601 (
            .O(N__49201),
            .I(N__48995));
    CascadeMux I__11600 (
            .O(N__49200),
            .I(N__48991));
    CascadeMux I__11599 (
            .O(N__49199),
            .I(N__48988));
    CascadeMux I__11598 (
            .O(N__49198),
            .I(N__48985));
    CascadeMux I__11597 (
            .O(N__49197),
            .I(N__48980));
    CascadeMux I__11596 (
            .O(N__49196),
            .I(N__48976));
    CascadeMux I__11595 (
            .O(N__49195),
            .I(N__48972));
    InMux I__11594 (
            .O(N__49192),
            .I(N__48955));
    InMux I__11593 (
            .O(N__49191),
            .I(N__48955));
    InMux I__11592 (
            .O(N__49188),
            .I(N__48955));
    InMux I__11591 (
            .O(N__49187),
            .I(N__48955));
    InMux I__11590 (
            .O(N__49184),
            .I(N__48955));
    InMux I__11589 (
            .O(N__49183),
            .I(N__48955));
    InMux I__11588 (
            .O(N__49180),
            .I(N__48955));
    InMux I__11587 (
            .O(N__49179),
            .I(N__48955));
    InMux I__11586 (
            .O(N__49178),
            .I(N__48942));
    InMux I__11585 (
            .O(N__49175),
            .I(N__48942));
    InMux I__11584 (
            .O(N__49174),
            .I(N__48942));
    InMux I__11583 (
            .O(N__49171),
            .I(N__48942));
    InMux I__11582 (
            .O(N__49170),
            .I(N__48942));
    InMux I__11581 (
            .O(N__49167),
            .I(N__48942));
    Span4Mux_h I__11580 (
            .O(N__49164),
            .I(N__48939));
    Sp12to4 I__11579 (
            .O(N__49159),
            .I(N__48936));
    Span4Mux_h I__11578 (
            .O(N__49154),
            .I(N__48931));
    LocalMux I__11577 (
            .O(N__49137),
            .I(N__48931));
    LocalMux I__11576 (
            .O(N__49128),
            .I(N__48926));
    LocalMux I__11575 (
            .O(N__49123),
            .I(N__48926));
    InMux I__11574 (
            .O(N__49120),
            .I(N__48917));
    InMux I__11573 (
            .O(N__49117),
            .I(N__48917));
    InMux I__11572 (
            .O(N__49114),
            .I(N__48917));
    InMux I__11571 (
            .O(N__49111),
            .I(N__48917));
    InMux I__11570 (
            .O(N__49110),
            .I(N__48912));
    InMux I__11569 (
            .O(N__49107),
            .I(N__48912));
    InMux I__11568 (
            .O(N__49106),
            .I(N__48903));
    InMux I__11567 (
            .O(N__49105),
            .I(N__48903));
    InMux I__11566 (
            .O(N__49104),
            .I(N__48903));
    InMux I__11565 (
            .O(N__49103),
            .I(N__48903));
    InMux I__11564 (
            .O(N__49100),
            .I(N__48900));
    InMux I__11563 (
            .O(N__49099),
            .I(N__48883));
    InMux I__11562 (
            .O(N__49096),
            .I(N__48883));
    InMux I__11561 (
            .O(N__49095),
            .I(N__48883));
    InMux I__11560 (
            .O(N__49092),
            .I(N__48883));
    InMux I__11559 (
            .O(N__49091),
            .I(N__48883));
    InMux I__11558 (
            .O(N__49088),
            .I(N__48883));
    InMux I__11557 (
            .O(N__49087),
            .I(N__48883));
    InMux I__11556 (
            .O(N__49084),
            .I(N__48883));
    InMux I__11555 (
            .O(N__49081),
            .I(N__48866));
    InMux I__11554 (
            .O(N__49080),
            .I(N__48866));
    InMux I__11553 (
            .O(N__49077),
            .I(N__48866));
    InMux I__11552 (
            .O(N__49076),
            .I(N__48866));
    InMux I__11551 (
            .O(N__49073),
            .I(N__48866));
    InMux I__11550 (
            .O(N__49072),
            .I(N__48866));
    InMux I__11549 (
            .O(N__49069),
            .I(N__48866));
    InMux I__11548 (
            .O(N__49068),
            .I(N__48866));
    Span4Mux_v I__11547 (
            .O(N__49065),
            .I(N__48849));
    LocalMux I__11546 (
            .O(N__49060),
            .I(N__48849));
    LocalMux I__11545 (
            .O(N__49055),
            .I(N__48849));
    LocalMux I__11544 (
            .O(N__49040),
            .I(N__48849));
    Span4Mux_h I__11543 (
            .O(N__49035),
            .I(N__48849));
    Span4Mux_h I__11542 (
            .O(N__49032),
            .I(N__48849));
    LocalMux I__11541 (
            .O(N__49021),
            .I(N__48849));
    LocalMux I__11540 (
            .O(N__49004),
            .I(N__48849));
    InMux I__11539 (
            .O(N__49001),
            .I(N__48840));
    InMux I__11538 (
            .O(N__48998),
            .I(N__48840));
    InMux I__11537 (
            .O(N__48995),
            .I(N__48840));
    InMux I__11536 (
            .O(N__48994),
            .I(N__48840));
    InMux I__11535 (
            .O(N__48991),
            .I(N__48831));
    InMux I__11534 (
            .O(N__48988),
            .I(N__48831));
    InMux I__11533 (
            .O(N__48985),
            .I(N__48831));
    InMux I__11532 (
            .O(N__48984),
            .I(N__48831));
    InMux I__11531 (
            .O(N__48983),
            .I(N__48818));
    InMux I__11530 (
            .O(N__48980),
            .I(N__48818));
    InMux I__11529 (
            .O(N__48979),
            .I(N__48818));
    InMux I__11528 (
            .O(N__48976),
            .I(N__48818));
    InMux I__11527 (
            .O(N__48975),
            .I(N__48818));
    InMux I__11526 (
            .O(N__48972),
            .I(N__48818));
    LocalMux I__11525 (
            .O(N__48955),
            .I(N__48813));
    LocalMux I__11524 (
            .O(N__48942),
            .I(N__48813));
    Odrv4 I__11523 (
            .O(N__48939),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__11522 (
            .O(N__48936),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11521 (
            .O(N__48931),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11520 (
            .O(N__48926),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11519 (
            .O(N__48917),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11518 (
            .O(N__48912),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11517 (
            .O(N__48903),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11516 (
            .O(N__48900),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11515 (
            .O(N__48883),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11514 (
            .O(N__48866),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11513 (
            .O(N__48849),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11512 (
            .O(N__48840),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11511 (
            .O(N__48831),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11510 (
            .O(N__48818),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11509 (
            .O(N__48813),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__11508 (
            .O(N__48782),
            .I(N__48779));
    LocalMux I__11507 (
            .O(N__48779),
            .I(N__48776));
    Span4Mux_h I__11506 (
            .O(N__48776),
            .I(N__48773));
    Odrv4 I__11505 (
            .O(N__48773),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__11504 (
            .O(N__48770),
            .I(N__48765));
    InMux I__11503 (
            .O(N__48769),
            .I(N__48760));
    InMux I__11502 (
            .O(N__48768),
            .I(N__48760));
    LocalMux I__11501 (
            .O(N__48765),
            .I(N__48755));
    LocalMux I__11500 (
            .O(N__48760),
            .I(N__48755));
    Span4Mux_h I__11499 (
            .O(N__48755),
            .I(N__48751));
    InMux I__11498 (
            .O(N__48754),
            .I(N__48748));
    Odrv4 I__11497 (
            .O(N__48751),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__11496 (
            .O(N__48748),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__11495 (
            .O(N__48743),
            .I(N__48734));
    InMux I__11494 (
            .O(N__48742),
            .I(N__48734));
    InMux I__11493 (
            .O(N__48741),
            .I(N__48734));
    LocalMux I__11492 (
            .O(N__48734),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__11491 (
            .O(N__48731),
            .I(N__48728));
    LocalMux I__11490 (
            .O(N__48728),
            .I(N__48725));
    Odrv12 I__11489 (
            .O(N__48725),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__11488 (
            .O(N__48722),
            .I(N__48718));
    InMux I__11487 (
            .O(N__48721),
            .I(N__48715));
    LocalMux I__11486 (
            .O(N__48718),
            .I(N__48712));
    LocalMux I__11485 (
            .O(N__48715),
            .I(N__48709));
    Span4Mux_h I__11484 (
            .O(N__48712),
            .I(N__48706));
    Span4Mux_h I__11483 (
            .O(N__48709),
            .I(N__48702));
    Span4Mux_v I__11482 (
            .O(N__48706),
            .I(N__48699));
    InMux I__11481 (
            .O(N__48705),
            .I(N__48696));
    Odrv4 I__11480 (
            .O(N__48702),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__11479 (
            .O(N__48699),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    LocalMux I__11478 (
            .O(N__48696),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__11477 (
            .O(N__48689),
            .I(N__48680));
    InMux I__11476 (
            .O(N__48688),
            .I(N__48680));
    InMux I__11475 (
            .O(N__48687),
            .I(N__48677));
    InMux I__11474 (
            .O(N__48686),
            .I(N__48662));
    CascadeMux I__11473 (
            .O(N__48685),
            .I(N__48659));
    LocalMux I__11472 (
            .O(N__48680),
            .I(N__48653));
    LocalMux I__11471 (
            .O(N__48677),
            .I(N__48653));
    InMux I__11470 (
            .O(N__48676),
            .I(N__48640));
    InMux I__11469 (
            .O(N__48675),
            .I(N__48640));
    InMux I__11468 (
            .O(N__48674),
            .I(N__48640));
    InMux I__11467 (
            .O(N__48673),
            .I(N__48640));
    InMux I__11466 (
            .O(N__48672),
            .I(N__48640));
    InMux I__11465 (
            .O(N__48671),
            .I(N__48640));
    InMux I__11464 (
            .O(N__48670),
            .I(N__48635));
    InMux I__11463 (
            .O(N__48669),
            .I(N__48635));
    InMux I__11462 (
            .O(N__48668),
            .I(N__48630));
    InMux I__11461 (
            .O(N__48667),
            .I(N__48630));
    InMux I__11460 (
            .O(N__48666),
            .I(N__48625));
    InMux I__11459 (
            .O(N__48665),
            .I(N__48625));
    LocalMux I__11458 (
            .O(N__48662),
            .I(N__48622));
    InMux I__11457 (
            .O(N__48659),
            .I(N__48617));
    InMux I__11456 (
            .O(N__48658),
            .I(N__48617));
    Span4Mux_v I__11455 (
            .O(N__48653),
            .I(N__48614));
    LocalMux I__11454 (
            .O(N__48640),
            .I(N__48609));
    LocalMux I__11453 (
            .O(N__48635),
            .I(N__48609));
    LocalMux I__11452 (
            .O(N__48630),
            .I(N__48598));
    LocalMux I__11451 (
            .O(N__48625),
            .I(N__48598));
    Span4Mux_h I__11450 (
            .O(N__48622),
            .I(N__48595));
    LocalMux I__11449 (
            .O(N__48617),
            .I(N__48588));
    Span4Mux_h I__11448 (
            .O(N__48614),
            .I(N__48588));
    Span4Mux_v I__11447 (
            .O(N__48609),
            .I(N__48588));
    InMux I__11446 (
            .O(N__48608),
            .I(N__48579));
    InMux I__11445 (
            .O(N__48607),
            .I(N__48579));
    InMux I__11444 (
            .O(N__48606),
            .I(N__48579));
    InMux I__11443 (
            .O(N__48605),
            .I(N__48579));
    InMux I__11442 (
            .O(N__48604),
            .I(N__48576));
    InMux I__11441 (
            .O(N__48603),
            .I(N__48572));
    Span4Mux_v I__11440 (
            .O(N__48598),
            .I(N__48569));
    Span4Mux_v I__11439 (
            .O(N__48595),
            .I(N__48566));
    Sp12to4 I__11438 (
            .O(N__48588),
            .I(N__48559));
    LocalMux I__11437 (
            .O(N__48579),
            .I(N__48559));
    LocalMux I__11436 (
            .O(N__48576),
            .I(N__48559));
    InMux I__11435 (
            .O(N__48575),
            .I(N__48556));
    LocalMux I__11434 (
            .O(N__48572),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__11433 (
            .O(N__48569),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__11432 (
            .O(N__48566),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv12 I__11431 (
            .O(N__48559),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__11430 (
            .O(N__48556),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__11429 (
            .O(N__48545),
            .I(N__48541));
    InMux I__11428 (
            .O(N__48544),
            .I(N__48538));
    InMux I__11427 (
            .O(N__48541),
            .I(N__48535));
    LocalMux I__11426 (
            .O(N__48538),
            .I(N__48532));
    LocalMux I__11425 (
            .O(N__48535),
            .I(N__48528));
    Span12Mux_s10_h I__11424 (
            .O(N__48532),
            .I(N__48525));
    InMux I__11423 (
            .O(N__48531),
            .I(N__48522));
    Span4Mux_v I__11422 (
            .O(N__48528),
            .I(N__48519));
    Odrv12 I__11421 (
            .O(N__48525),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__11420 (
            .O(N__48522),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__11419 (
            .O(N__48519),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__11418 (
            .O(N__48512),
            .I(N__48509));
    LocalMux I__11417 (
            .O(N__48509),
            .I(N__48505));
    InMux I__11416 (
            .O(N__48508),
            .I(N__48502));
    Span4Mux_h I__11415 (
            .O(N__48505),
            .I(N__48497));
    LocalMux I__11414 (
            .O(N__48502),
            .I(N__48497));
    Span4Mux_v I__11413 (
            .O(N__48497),
            .I(N__48492));
    InMux I__11412 (
            .O(N__48496),
            .I(N__48487));
    InMux I__11411 (
            .O(N__48495),
            .I(N__48487));
    Odrv4 I__11410 (
            .O(N__48492),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__11409 (
            .O(N__48487),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    ClkMux I__11408 (
            .O(N__48482),
            .I(N__48020));
    ClkMux I__11407 (
            .O(N__48481),
            .I(N__48020));
    ClkMux I__11406 (
            .O(N__48480),
            .I(N__48020));
    ClkMux I__11405 (
            .O(N__48479),
            .I(N__48020));
    ClkMux I__11404 (
            .O(N__48478),
            .I(N__48020));
    ClkMux I__11403 (
            .O(N__48477),
            .I(N__48020));
    ClkMux I__11402 (
            .O(N__48476),
            .I(N__48020));
    ClkMux I__11401 (
            .O(N__48475),
            .I(N__48020));
    ClkMux I__11400 (
            .O(N__48474),
            .I(N__48020));
    ClkMux I__11399 (
            .O(N__48473),
            .I(N__48020));
    ClkMux I__11398 (
            .O(N__48472),
            .I(N__48020));
    ClkMux I__11397 (
            .O(N__48471),
            .I(N__48020));
    ClkMux I__11396 (
            .O(N__48470),
            .I(N__48020));
    ClkMux I__11395 (
            .O(N__48469),
            .I(N__48020));
    ClkMux I__11394 (
            .O(N__48468),
            .I(N__48020));
    ClkMux I__11393 (
            .O(N__48467),
            .I(N__48020));
    ClkMux I__11392 (
            .O(N__48466),
            .I(N__48020));
    ClkMux I__11391 (
            .O(N__48465),
            .I(N__48020));
    ClkMux I__11390 (
            .O(N__48464),
            .I(N__48020));
    ClkMux I__11389 (
            .O(N__48463),
            .I(N__48020));
    ClkMux I__11388 (
            .O(N__48462),
            .I(N__48020));
    ClkMux I__11387 (
            .O(N__48461),
            .I(N__48020));
    ClkMux I__11386 (
            .O(N__48460),
            .I(N__48020));
    ClkMux I__11385 (
            .O(N__48459),
            .I(N__48020));
    ClkMux I__11384 (
            .O(N__48458),
            .I(N__48020));
    ClkMux I__11383 (
            .O(N__48457),
            .I(N__48020));
    ClkMux I__11382 (
            .O(N__48456),
            .I(N__48020));
    ClkMux I__11381 (
            .O(N__48455),
            .I(N__48020));
    ClkMux I__11380 (
            .O(N__48454),
            .I(N__48020));
    ClkMux I__11379 (
            .O(N__48453),
            .I(N__48020));
    ClkMux I__11378 (
            .O(N__48452),
            .I(N__48020));
    ClkMux I__11377 (
            .O(N__48451),
            .I(N__48020));
    ClkMux I__11376 (
            .O(N__48450),
            .I(N__48020));
    ClkMux I__11375 (
            .O(N__48449),
            .I(N__48020));
    ClkMux I__11374 (
            .O(N__48448),
            .I(N__48020));
    ClkMux I__11373 (
            .O(N__48447),
            .I(N__48020));
    ClkMux I__11372 (
            .O(N__48446),
            .I(N__48020));
    ClkMux I__11371 (
            .O(N__48445),
            .I(N__48020));
    ClkMux I__11370 (
            .O(N__48444),
            .I(N__48020));
    ClkMux I__11369 (
            .O(N__48443),
            .I(N__48020));
    ClkMux I__11368 (
            .O(N__48442),
            .I(N__48020));
    ClkMux I__11367 (
            .O(N__48441),
            .I(N__48020));
    ClkMux I__11366 (
            .O(N__48440),
            .I(N__48020));
    ClkMux I__11365 (
            .O(N__48439),
            .I(N__48020));
    ClkMux I__11364 (
            .O(N__48438),
            .I(N__48020));
    ClkMux I__11363 (
            .O(N__48437),
            .I(N__48020));
    ClkMux I__11362 (
            .O(N__48436),
            .I(N__48020));
    ClkMux I__11361 (
            .O(N__48435),
            .I(N__48020));
    ClkMux I__11360 (
            .O(N__48434),
            .I(N__48020));
    ClkMux I__11359 (
            .O(N__48433),
            .I(N__48020));
    ClkMux I__11358 (
            .O(N__48432),
            .I(N__48020));
    ClkMux I__11357 (
            .O(N__48431),
            .I(N__48020));
    ClkMux I__11356 (
            .O(N__48430),
            .I(N__48020));
    ClkMux I__11355 (
            .O(N__48429),
            .I(N__48020));
    ClkMux I__11354 (
            .O(N__48428),
            .I(N__48020));
    ClkMux I__11353 (
            .O(N__48427),
            .I(N__48020));
    ClkMux I__11352 (
            .O(N__48426),
            .I(N__48020));
    ClkMux I__11351 (
            .O(N__48425),
            .I(N__48020));
    ClkMux I__11350 (
            .O(N__48424),
            .I(N__48020));
    ClkMux I__11349 (
            .O(N__48423),
            .I(N__48020));
    ClkMux I__11348 (
            .O(N__48422),
            .I(N__48020));
    ClkMux I__11347 (
            .O(N__48421),
            .I(N__48020));
    ClkMux I__11346 (
            .O(N__48420),
            .I(N__48020));
    ClkMux I__11345 (
            .O(N__48419),
            .I(N__48020));
    ClkMux I__11344 (
            .O(N__48418),
            .I(N__48020));
    ClkMux I__11343 (
            .O(N__48417),
            .I(N__48020));
    ClkMux I__11342 (
            .O(N__48416),
            .I(N__48020));
    ClkMux I__11341 (
            .O(N__48415),
            .I(N__48020));
    ClkMux I__11340 (
            .O(N__48414),
            .I(N__48020));
    ClkMux I__11339 (
            .O(N__48413),
            .I(N__48020));
    ClkMux I__11338 (
            .O(N__48412),
            .I(N__48020));
    ClkMux I__11337 (
            .O(N__48411),
            .I(N__48020));
    ClkMux I__11336 (
            .O(N__48410),
            .I(N__48020));
    ClkMux I__11335 (
            .O(N__48409),
            .I(N__48020));
    ClkMux I__11334 (
            .O(N__48408),
            .I(N__48020));
    ClkMux I__11333 (
            .O(N__48407),
            .I(N__48020));
    ClkMux I__11332 (
            .O(N__48406),
            .I(N__48020));
    ClkMux I__11331 (
            .O(N__48405),
            .I(N__48020));
    ClkMux I__11330 (
            .O(N__48404),
            .I(N__48020));
    ClkMux I__11329 (
            .O(N__48403),
            .I(N__48020));
    ClkMux I__11328 (
            .O(N__48402),
            .I(N__48020));
    ClkMux I__11327 (
            .O(N__48401),
            .I(N__48020));
    ClkMux I__11326 (
            .O(N__48400),
            .I(N__48020));
    ClkMux I__11325 (
            .O(N__48399),
            .I(N__48020));
    ClkMux I__11324 (
            .O(N__48398),
            .I(N__48020));
    ClkMux I__11323 (
            .O(N__48397),
            .I(N__48020));
    ClkMux I__11322 (
            .O(N__48396),
            .I(N__48020));
    ClkMux I__11321 (
            .O(N__48395),
            .I(N__48020));
    ClkMux I__11320 (
            .O(N__48394),
            .I(N__48020));
    ClkMux I__11319 (
            .O(N__48393),
            .I(N__48020));
    ClkMux I__11318 (
            .O(N__48392),
            .I(N__48020));
    ClkMux I__11317 (
            .O(N__48391),
            .I(N__48020));
    ClkMux I__11316 (
            .O(N__48390),
            .I(N__48020));
    ClkMux I__11315 (
            .O(N__48389),
            .I(N__48020));
    ClkMux I__11314 (
            .O(N__48388),
            .I(N__48020));
    ClkMux I__11313 (
            .O(N__48387),
            .I(N__48020));
    ClkMux I__11312 (
            .O(N__48386),
            .I(N__48020));
    ClkMux I__11311 (
            .O(N__48385),
            .I(N__48020));
    ClkMux I__11310 (
            .O(N__48384),
            .I(N__48020));
    ClkMux I__11309 (
            .O(N__48383),
            .I(N__48020));
    ClkMux I__11308 (
            .O(N__48382),
            .I(N__48020));
    ClkMux I__11307 (
            .O(N__48381),
            .I(N__48020));
    ClkMux I__11306 (
            .O(N__48380),
            .I(N__48020));
    ClkMux I__11305 (
            .O(N__48379),
            .I(N__48020));
    ClkMux I__11304 (
            .O(N__48378),
            .I(N__48020));
    ClkMux I__11303 (
            .O(N__48377),
            .I(N__48020));
    ClkMux I__11302 (
            .O(N__48376),
            .I(N__48020));
    ClkMux I__11301 (
            .O(N__48375),
            .I(N__48020));
    ClkMux I__11300 (
            .O(N__48374),
            .I(N__48020));
    ClkMux I__11299 (
            .O(N__48373),
            .I(N__48020));
    ClkMux I__11298 (
            .O(N__48372),
            .I(N__48020));
    ClkMux I__11297 (
            .O(N__48371),
            .I(N__48020));
    ClkMux I__11296 (
            .O(N__48370),
            .I(N__48020));
    ClkMux I__11295 (
            .O(N__48369),
            .I(N__48020));
    ClkMux I__11294 (
            .O(N__48368),
            .I(N__48020));
    ClkMux I__11293 (
            .O(N__48367),
            .I(N__48020));
    ClkMux I__11292 (
            .O(N__48366),
            .I(N__48020));
    ClkMux I__11291 (
            .O(N__48365),
            .I(N__48020));
    ClkMux I__11290 (
            .O(N__48364),
            .I(N__48020));
    ClkMux I__11289 (
            .O(N__48363),
            .I(N__48020));
    ClkMux I__11288 (
            .O(N__48362),
            .I(N__48020));
    ClkMux I__11287 (
            .O(N__48361),
            .I(N__48020));
    ClkMux I__11286 (
            .O(N__48360),
            .I(N__48020));
    ClkMux I__11285 (
            .O(N__48359),
            .I(N__48020));
    ClkMux I__11284 (
            .O(N__48358),
            .I(N__48020));
    ClkMux I__11283 (
            .O(N__48357),
            .I(N__48020));
    ClkMux I__11282 (
            .O(N__48356),
            .I(N__48020));
    ClkMux I__11281 (
            .O(N__48355),
            .I(N__48020));
    ClkMux I__11280 (
            .O(N__48354),
            .I(N__48020));
    ClkMux I__11279 (
            .O(N__48353),
            .I(N__48020));
    ClkMux I__11278 (
            .O(N__48352),
            .I(N__48020));
    ClkMux I__11277 (
            .O(N__48351),
            .I(N__48020));
    ClkMux I__11276 (
            .O(N__48350),
            .I(N__48020));
    ClkMux I__11275 (
            .O(N__48349),
            .I(N__48020));
    ClkMux I__11274 (
            .O(N__48348),
            .I(N__48020));
    ClkMux I__11273 (
            .O(N__48347),
            .I(N__48020));
    ClkMux I__11272 (
            .O(N__48346),
            .I(N__48020));
    ClkMux I__11271 (
            .O(N__48345),
            .I(N__48020));
    ClkMux I__11270 (
            .O(N__48344),
            .I(N__48020));
    ClkMux I__11269 (
            .O(N__48343),
            .I(N__48020));
    ClkMux I__11268 (
            .O(N__48342),
            .I(N__48020));
    ClkMux I__11267 (
            .O(N__48341),
            .I(N__48020));
    ClkMux I__11266 (
            .O(N__48340),
            .I(N__48020));
    ClkMux I__11265 (
            .O(N__48339),
            .I(N__48020));
    ClkMux I__11264 (
            .O(N__48338),
            .I(N__48020));
    ClkMux I__11263 (
            .O(N__48337),
            .I(N__48020));
    ClkMux I__11262 (
            .O(N__48336),
            .I(N__48020));
    ClkMux I__11261 (
            .O(N__48335),
            .I(N__48020));
    ClkMux I__11260 (
            .O(N__48334),
            .I(N__48020));
    ClkMux I__11259 (
            .O(N__48333),
            .I(N__48020));
    ClkMux I__11258 (
            .O(N__48332),
            .I(N__48020));
    ClkMux I__11257 (
            .O(N__48331),
            .I(N__48020));
    ClkMux I__11256 (
            .O(N__48330),
            .I(N__48020));
    ClkMux I__11255 (
            .O(N__48329),
            .I(N__48020));
    GlobalMux I__11254 (
            .O(N__48020),
            .I(clk_100mhz_0));
    CEMux I__11253 (
            .O(N__48017),
            .I(N__48013));
    CEMux I__11252 (
            .O(N__48016),
            .I(N__48009));
    LocalMux I__11251 (
            .O(N__48013),
            .I(N__48005));
    CEMux I__11250 (
            .O(N__48012),
            .I(N__48002));
    LocalMux I__11249 (
            .O(N__48009),
            .I(N__47999));
    CEMux I__11248 (
            .O(N__48008),
            .I(N__47996));
    Span4Mux_v I__11247 (
            .O(N__48005),
            .I(N__47989));
    LocalMux I__11246 (
            .O(N__48002),
            .I(N__47989));
    Span4Mux_h I__11245 (
            .O(N__47999),
            .I(N__47982));
    LocalMux I__11244 (
            .O(N__47996),
            .I(N__47982));
    CEMux I__11243 (
            .O(N__47995),
            .I(N__47979));
    CEMux I__11242 (
            .O(N__47994),
            .I(N__47976));
    Span4Mux_v I__11241 (
            .O(N__47989),
            .I(N__47973));
    CEMux I__11240 (
            .O(N__47988),
            .I(N__47970));
    CEMux I__11239 (
            .O(N__47987),
            .I(N__47967));
    Span4Mux_h I__11238 (
            .O(N__47982),
            .I(N__47960));
    LocalMux I__11237 (
            .O(N__47979),
            .I(N__47960));
    LocalMux I__11236 (
            .O(N__47976),
            .I(N__47960));
    Span4Mux_h I__11235 (
            .O(N__47973),
            .I(N__47955));
    LocalMux I__11234 (
            .O(N__47970),
            .I(N__47955));
    LocalMux I__11233 (
            .O(N__47967),
            .I(N__47951));
    Span4Mux_v I__11232 (
            .O(N__47960),
            .I(N__47948));
    Span4Mux_h I__11231 (
            .O(N__47955),
            .I(N__47945));
    CEMux I__11230 (
            .O(N__47954),
            .I(N__47942));
    Span4Mux_v I__11229 (
            .O(N__47951),
            .I(N__47937));
    Span4Mux_h I__11228 (
            .O(N__47948),
            .I(N__47937));
    Span4Mux_v I__11227 (
            .O(N__47945),
            .I(N__47932));
    LocalMux I__11226 (
            .O(N__47942),
            .I(N__47932));
    Odrv4 I__11225 (
            .O(N__47937),
            .I(\current_shift_inst.timer_s1.N_180_i_g ));
    Odrv4 I__11224 (
            .O(N__47932),
            .I(\current_shift_inst.timer_s1.N_180_i_g ));
    CascadeMux I__11223 (
            .O(N__47927),
            .I(N__47919));
    CascadeMux I__11222 (
            .O(N__47926),
            .I(N__47915));
    InMux I__11221 (
            .O(N__47925),
            .I(N__47912));
    InMux I__11220 (
            .O(N__47924),
            .I(N__47909));
    InMux I__11219 (
            .O(N__47923),
            .I(N__47906));
    InMux I__11218 (
            .O(N__47922),
            .I(N__47903));
    InMux I__11217 (
            .O(N__47919),
            .I(N__47900));
    InMux I__11216 (
            .O(N__47918),
            .I(N__47897));
    InMux I__11215 (
            .O(N__47915),
            .I(N__47894));
    LocalMux I__11214 (
            .O(N__47912),
            .I(N__47891));
    LocalMux I__11213 (
            .O(N__47909),
            .I(N__47888));
    LocalMux I__11212 (
            .O(N__47906),
            .I(N__47885));
    LocalMux I__11211 (
            .O(N__47903),
            .I(N__47844));
    LocalMux I__11210 (
            .O(N__47900),
            .I(N__47781));
    LocalMux I__11209 (
            .O(N__47897),
            .I(N__47762));
    LocalMux I__11208 (
            .O(N__47894),
            .I(N__47743));
    Glb2LocalMux I__11207 (
            .O(N__47891),
            .I(N__47444));
    Glb2LocalMux I__11206 (
            .O(N__47888),
            .I(N__47444));
    Glb2LocalMux I__11205 (
            .O(N__47885),
            .I(N__47444));
    SRMux I__11204 (
            .O(N__47884),
            .I(N__47444));
    SRMux I__11203 (
            .O(N__47883),
            .I(N__47444));
    SRMux I__11202 (
            .O(N__47882),
            .I(N__47444));
    SRMux I__11201 (
            .O(N__47881),
            .I(N__47444));
    SRMux I__11200 (
            .O(N__47880),
            .I(N__47444));
    SRMux I__11199 (
            .O(N__47879),
            .I(N__47444));
    SRMux I__11198 (
            .O(N__47878),
            .I(N__47444));
    SRMux I__11197 (
            .O(N__47877),
            .I(N__47444));
    SRMux I__11196 (
            .O(N__47876),
            .I(N__47444));
    SRMux I__11195 (
            .O(N__47875),
            .I(N__47444));
    SRMux I__11194 (
            .O(N__47874),
            .I(N__47444));
    SRMux I__11193 (
            .O(N__47873),
            .I(N__47444));
    SRMux I__11192 (
            .O(N__47872),
            .I(N__47444));
    SRMux I__11191 (
            .O(N__47871),
            .I(N__47444));
    SRMux I__11190 (
            .O(N__47870),
            .I(N__47444));
    SRMux I__11189 (
            .O(N__47869),
            .I(N__47444));
    SRMux I__11188 (
            .O(N__47868),
            .I(N__47444));
    SRMux I__11187 (
            .O(N__47867),
            .I(N__47444));
    SRMux I__11186 (
            .O(N__47866),
            .I(N__47444));
    SRMux I__11185 (
            .O(N__47865),
            .I(N__47444));
    SRMux I__11184 (
            .O(N__47864),
            .I(N__47444));
    SRMux I__11183 (
            .O(N__47863),
            .I(N__47444));
    SRMux I__11182 (
            .O(N__47862),
            .I(N__47444));
    SRMux I__11181 (
            .O(N__47861),
            .I(N__47444));
    SRMux I__11180 (
            .O(N__47860),
            .I(N__47444));
    SRMux I__11179 (
            .O(N__47859),
            .I(N__47444));
    SRMux I__11178 (
            .O(N__47858),
            .I(N__47444));
    SRMux I__11177 (
            .O(N__47857),
            .I(N__47444));
    SRMux I__11176 (
            .O(N__47856),
            .I(N__47444));
    SRMux I__11175 (
            .O(N__47855),
            .I(N__47444));
    SRMux I__11174 (
            .O(N__47854),
            .I(N__47444));
    SRMux I__11173 (
            .O(N__47853),
            .I(N__47444));
    SRMux I__11172 (
            .O(N__47852),
            .I(N__47444));
    SRMux I__11171 (
            .O(N__47851),
            .I(N__47444));
    SRMux I__11170 (
            .O(N__47850),
            .I(N__47444));
    SRMux I__11169 (
            .O(N__47849),
            .I(N__47444));
    SRMux I__11168 (
            .O(N__47848),
            .I(N__47444));
    SRMux I__11167 (
            .O(N__47847),
            .I(N__47444));
    Glb2LocalMux I__11166 (
            .O(N__47844),
            .I(N__47444));
    SRMux I__11165 (
            .O(N__47843),
            .I(N__47444));
    SRMux I__11164 (
            .O(N__47842),
            .I(N__47444));
    SRMux I__11163 (
            .O(N__47841),
            .I(N__47444));
    SRMux I__11162 (
            .O(N__47840),
            .I(N__47444));
    SRMux I__11161 (
            .O(N__47839),
            .I(N__47444));
    SRMux I__11160 (
            .O(N__47838),
            .I(N__47444));
    SRMux I__11159 (
            .O(N__47837),
            .I(N__47444));
    SRMux I__11158 (
            .O(N__47836),
            .I(N__47444));
    SRMux I__11157 (
            .O(N__47835),
            .I(N__47444));
    SRMux I__11156 (
            .O(N__47834),
            .I(N__47444));
    SRMux I__11155 (
            .O(N__47833),
            .I(N__47444));
    SRMux I__11154 (
            .O(N__47832),
            .I(N__47444));
    SRMux I__11153 (
            .O(N__47831),
            .I(N__47444));
    SRMux I__11152 (
            .O(N__47830),
            .I(N__47444));
    SRMux I__11151 (
            .O(N__47829),
            .I(N__47444));
    SRMux I__11150 (
            .O(N__47828),
            .I(N__47444));
    SRMux I__11149 (
            .O(N__47827),
            .I(N__47444));
    SRMux I__11148 (
            .O(N__47826),
            .I(N__47444));
    SRMux I__11147 (
            .O(N__47825),
            .I(N__47444));
    SRMux I__11146 (
            .O(N__47824),
            .I(N__47444));
    SRMux I__11145 (
            .O(N__47823),
            .I(N__47444));
    SRMux I__11144 (
            .O(N__47822),
            .I(N__47444));
    SRMux I__11143 (
            .O(N__47821),
            .I(N__47444));
    SRMux I__11142 (
            .O(N__47820),
            .I(N__47444));
    SRMux I__11141 (
            .O(N__47819),
            .I(N__47444));
    SRMux I__11140 (
            .O(N__47818),
            .I(N__47444));
    SRMux I__11139 (
            .O(N__47817),
            .I(N__47444));
    SRMux I__11138 (
            .O(N__47816),
            .I(N__47444));
    SRMux I__11137 (
            .O(N__47815),
            .I(N__47444));
    SRMux I__11136 (
            .O(N__47814),
            .I(N__47444));
    SRMux I__11135 (
            .O(N__47813),
            .I(N__47444));
    SRMux I__11134 (
            .O(N__47812),
            .I(N__47444));
    SRMux I__11133 (
            .O(N__47811),
            .I(N__47444));
    SRMux I__11132 (
            .O(N__47810),
            .I(N__47444));
    SRMux I__11131 (
            .O(N__47809),
            .I(N__47444));
    SRMux I__11130 (
            .O(N__47808),
            .I(N__47444));
    SRMux I__11129 (
            .O(N__47807),
            .I(N__47444));
    SRMux I__11128 (
            .O(N__47806),
            .I(N__47444));
    SRMux I__11127 (
            .O(N__47805),
            .I(N__47444));
    SRMux I__11126 (
            .O(N__47804),
            .I(N__47444));
    SRMux I__11125 (
            .O(N__47803),
            .I(N__47444));
    SRMux I__11124 (
            .O(N__47802),
            .I(N__47444));
    SRMux I__11123 (
            .O(N__47801),
            .I(N__47444));
    SRMux I__11122 (
            .O(N__47800),
            .I(N__47444));
    SRMux I__11121 (
            .O(N__47799),
            .I(N__47444));
    SRMux I__11120 (
            .O(N__47798),
            .I(N__47444));
    SRMux I__11119 (
            .O(N__47797),
            .I(N__47444));
    SRMux I__11118 (
            .O(N__47796),
            .I(N__47444));
    SRMux I__11117 (
            .O(N__47795),
            .I(N__47444));
    SRMux I__11116 (
            .O(N__47794),
            .I(N__47444));
    SRMux I__11115 (
            .O(N__47793),
            .I(N__47444));
    SRMux I__11114 (
            .O(N__47792),
            .I(N__47444));
    SRMux I__11113 (
            .O(N__47791),
            .I(N__47444));
    SRMux I__11112 (
            .O(N__47790),
            .I(N__47444));
    SRMux I__11111 (
            .O(N__47789),
            .I(N__47444));
    SRMux I__11110 (
            .O(N__47788),
            .I(N__47444));
    SRMux I__11109 (
            .O(N__47787),
            .I(N__47444));
    SRMux I__11108 (
            .O(N__47786),
            .I(N__47444));
    SRMux I__11107 (
            .O(N__47785),
            .I(N__47444));
    SRMux I__11106 (
            .O(N__47784),
            .I(N__47444));
    Glb2LocalMux I__11105 (
            .O(N__47781),
            .I(N__47444));
    SRMux I__11104 (
            .O(N__47780),
            .I(N__47444));
    SRMux I__11103 (
            .O(N__47779),
            .I(N__47444));
    SRMux I__11102 (
            .O(N__47778),
            .I(N__47444));
    SRMux I__11101 (
            .O(N__47777),
            .I(N__47444));
    SRMux I__11100 (
            .O(N__47776),
            .I(N__47444));
    SRMux I__11099 (
            .O(N__47775),
            .I(N__47444));
    SRMux I__11098 (
            .O(N__47774),
            .I(N__47444));
    SRMux I__11097 (
            .O(N__47773),
            .I(N__47444));
    SRMux I__11096 (
            .O(N__47772),
            .I(N__47444));
    SRMux I__11095 (
            .O(N__47771),
            .I(N__47444));
    SRMux I__11094 (
            .O(N__47770),
            .I(N__47444));
    SRMux I__11093 (
            .O(N__47769),
            .I(N__47444));
    SRMux I__11092 (
            .O(N__47768),
            .I(N__47444));
    SRMux I__11091 (
            .O(N__47767),
            .I(N__47444));
    SRMux I__11090 (
            .O(N__47766),
            .I(N__47444));
    SRMux I__11089 (
            .O(N__47765),
            .I(N__47444));
    Glb2LocalMux I__11088 (
            .O(N__47762),
            .I(N__47444));
    SRMux I__11087 (
            .O(N__47761),
            .I(N__47444));
    SRMux I__11086 (
            .O(N__47760),
            .I(N__47444));
    SRMux I__11085 (
            .O(N__47759),
            .I(N__47444));
    SRMux I__11084 (
            .O(N__47758),
            .I(N__47444));
    SRMux I__11083 (
            .O(N__47757),
            .I(N__47444));
    SRMux I__11082 (
            .O(N__47756),
            .I(N__47444));
    SRMux I__11081 (
            .O(N__47755),
            .I(N__47444));
    SRMux I__11080 (
            .O(N__47754),
            .I(N__47444));
    SRMux I__11079 (
            .O(N__47753),
            .I(N__47444));
    SRMux I__11078 (
            .O(N__47752),
            .I(N__47444));
    SRMux I__11077 (
            .O(N__47751),
            .I(N__47444));
    SRMux I__11076 (
            .O(N__47750),
            .I(N__47444));
    SRMux I__11075 (
            .O(N__47749),
            .I(N__47444));
    SRMux I__11074 (
            .O(N__47748),
            .I(N__47444));
    SRMux I__11073 (
            .O(N__47747),
            .I(N__47444));
    SRMux I__11072 (
            .O(N__47746),
            .I(N__47444));
    Glb2LocalMux I__11071 (
            .O(N__47743),
            .I(N__47444));
    SRMux I__11070 (
            .O(N__47742),
            .I(N__47444));
    SRMux I__11069 (
            .O(N__47741),
            .I(N__47444));
    SRMux I__11068 (
            .O(N__47740),
            .I(N__47444));
    SRMux I__11067 (
            .O(N__47739),
            .I(N__47444));
    SRMux I__11066 (
            .O(N__47738),
            .I(N__47444));
    SRMux I__11065 (
            .O(N__47737),
            .I(N__47444));
    SRMux I__11064 (
            .O(N__47736),
            .I(N__47444));
    SRMux I__11063 (
            .O(N__47735),
            .I(N__47444));
    GlobalMux I__11062 (
            .O(N__47444),
            .I(N__47441));
    gio2CtrlBuf I__11061 (
            .O(N__47441),
            .I(red_c_g));
    CascadeMux I__11060 (
            .O(N__47438),
            .I(N__47434));
    InMux I__11059 (
            .O(N__47437),
            .I(N__47431));
    InMux I__11058 (
            .O(N__47434),
            .I(N__47428));
    LocalMux I__11057 (
            .O(N__47431),
            .I(N__47423));
    LocalMux I__11056 (
            .O(N__47428),
            .I(N__47420));
    InMux I__11055 (
            .O(N__47427),
            .I(N__47417));
    InMux I__11054 (
            .O(N__47426),
            .I(N__47414));
    Span4Mux_h I__11053 (
            .O(N__47423),
            .I(N__47411));
    Span4Mux_v I__11052 (
            .O(N__47420),
            .I(N__47408));
    LocalMux I__11051 (
            .O(N__47417),
            .I(N__47403));
    LocalMux I__11050 (
            .O(N__47414),
            .I(N__47403));
    Span4Mux_v I__11049 (
            .O(N__47411),
            .I(N__47398));
    Span4Mux_v I__11048 (
            .O(N__47408),
            .I(N__47398));
    Span4Mux_h I__11047 (
            .O(N__47403),
            .I(N__47395));
    Odrv4 I__11046 (
            .O(N__47398),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__11045 (
            .O(N__47395),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__11044 (
            .O(N__47390),
            .I(N__47387));
    LocalMux I__11043 (
            .O(N__47387),
            .I(N__47382));
    InMux I__11042 (
            .O(N__47386),
            .I(N__47379));
    InMux I__11041 (
            .O(N__47385),
            .I(N__47376));
    Odrv4 I__11040 (
            .O(N__47382),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__11039 (
            .O(N__47379),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__11038 (
            .O(N__47376),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__11037 (
            .O(N__47369),
            .I(N__47366));
    LocalMux I__11036 (
            .O(N__47366),
            .I(N__47363));
    Span4Mux_v I__11035 (
            .O(N__47363),
            .I(N__47360));
    Odrv4 I__11034 (
            .O(N__47360),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__11033 (
            .O(N__47357),
            .I(N__47353));
    InMux I__11032 (
            .O(N__47356),
            .I(N__47350));
    LocalMux I__11031 (
            .O(N__47353),
            .I(N__47346));
    LocalMux I__11030 (
            .O(N__47350),
            .I(N__47343));
    InMux I__11029 (
            .O(N__47349),
            .I(N__47340));
    Span4Mux_v I__11028 (
            .O(N__47346),
            .I(N__47337));
    Span4Mux_v I__11027 (
            .O(N__47343),
            .I(N__47331));
    LocalMux I__11026 (
            .O(N__47340),
            .I(N__47331));
    Span4Mux_h I__11025 (
            .O(N__47337),
            .I(N__47328));
    InMux I__11024 (
            .O(N__47336),
            .I(N__47325));
    Odrv4 I__11023 (
            .O(N__47331),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__11022 (
            .O(N__47328),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__11021 (
            .O(N__47325),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    CascadeMux I__11020 (
            .O(N__47318),
            .I(N__47314));
    InMux I__11019 (
            .O(N__47317),
            .I(N__47310));
    InMux I__11018 (
            .O(N__47314),
            .I(N__47307));
    InMux I__11017 (
            .O(N__47313),
            .I(N__47304));
    LocalMux I__11016 (
            .O(N__47310),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__11015 (
            .O(N__47307),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__11014 (
            .O(N__47304),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__11013 (
            .O(N__47297),
            .I(N__47294));
    LocalMux I__11012 (
            .O(N__47294),
            .I(N__47291));
    Odrv4 I__11011 (
            .O(N__47291),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__11010 (
            .O(N__47288),
            .I(N__47283));
    InMux I__11009 (
            .O(N__47287),
            .I(N__47277));
    InMux I__11008 (
            .O(N__47286),
            .I(N__47277));
    LocalMux I__11007 (
            .O(N__47283),
            .I(N__47274));
    InMux I__11006 (
            .O(N__47282),
            .I(N__47271));
    LocalMux I__11005 (
            .O(N__47277),
            .I(N__47268));
    Span4Mux_h I__11004 (
            .O(N__47274),
            .I(N__47265));
    LocalMux I__11003 (
            .O(N__47271),
            .I(N__47260));
    Span4Mux_h I__11002 (
            .O(N__47268),
            .I(N__47260));
    Odrv4 I__11001 (
            .O(N__47265),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__11000 (
            .O(N__47260),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__10999 (
            .O(N__47255),
            .I(N__47250));
    InMux I__10998 (
            .O(N__47254),
            .I(N__47247));
    InMux I__10997 (
            .O(N__47253),
            .I(N__47244));
    LocalMux I__10996 (
            .O(N__47250),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__10995 (
            .O(N__47247),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__10994 (
            .O(N__47244),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__10993 (
            .O(N__47237),
            .I(N__47234));
    LocalMux I__10992 (
            .O(N__47234),
            .I(N__47231));
    Odrv12 I__10991 (
            .O(N__47231),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__10990 (
            .O(N__47228),
            .I(N__47224));
    InMux I__10989 (
            .O(N__47227),
            .I(N__47220));
    InMux I__10988 (
            .O(N__47224),
            .I(N__47217));
    InMux I__10987 (
            .O(N__47223),
            .I(N__47214));
    LocalMux I__10986 (
            .O(N__47220),
            .I(N__47211));
    LocalMux I__10985 (
            .O(N__47217),
            .I(N__47206));
    LocalMux I__10984 (
            .O(N__47214),
            .I(N__47206));
    Span4Mux_h I__10983 (
            .O(N__47211),
            .I(N__47202));
    Span4Mux_v I__10982 (
            .O(N__47206),
            .I(N__47199));
    InMux I__10981 (
            .O(N__47205),
            .I(N__47196));
    Span4Mux_v I__10980 (
            .O(N__47202),
            .I(N__47189));
    Span4Mux_v I__10979 (
            .O(N__47199),
            .I(N__47189));
    LocalMux I__10978 (
            .O(N__47196),
            .I(N__47189));
    Odrv4 I__10977 (
            .O(N__47189),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__10976 (
            .O(N__47186),
            .I(N__47181));
    InMux I__10975 (
            .O(N__47185),
            .I(N__47178));
    InMux I__10974 (
            .O(N__47184),
            .I(N__47175));
    LocalMux I__10973 (
            .O(N__47181),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__10972 (
            .O(N__47178),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__10971 (
            .O(N__47175),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__10970 (
            .O(N__47168),
            .I(N__47165));
    LocalMux I__10969 (
            .O(N__47165),
            .I(N__47162));
    Odrv4 I__10968 (
            .O(N__47162),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__10967 (
            .O(N__47159),
            .I(N__47155));
    InMux I__10966 (
            .O(N__47158),
            .I(N__47152));
    LocalMux I__10965 (
            .O(N__47155),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    LocalMux I__10964 (
            .O(N__47152),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__10963 (
            .O(N__47147),
            .I(N__47144));
    LocalMux I__10962 (
            .O(N__47144),
            .I(N__47141));
    Odrv4 I__10961 (
            .O(N__47141),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__10960 (
            .O(N__47138),
            .I(N__47133));
    InMux I__10959 (
            .O(N__47137),
            .I(N__47130));
    InMux I__10958 (
            .O(N__47136),
            .I(N__47127));
    LocalMux I__10957 (
            .O(N__47133),
            .I(N__47124));
    LocalMux I__10956 (
            .O(N__47130),
            .I(N__47121));
    LocalMux I__10955 (
            .O(N__47127),
            .I(N__47116));
    Span4Mux_v I__10954 (
            .O(N__47124),
            .I(N__47116));
    Span4Mux_v I__10953 (
            .O(N__47121),
            .I(N__47110));
    Span4Mux_h I__10952 (
            .O(N__47116),
            .I(N__47110));
    InMux I__10951 (
            .O(N__47115),
            .I(N__47107));
    Odrv4 I__10950 (
            .O(N__47110),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__10949 (
            .O(N__47107),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__10948 (
            .O(N__47102),
            .I(N__47099));
    LocalMux I__10947 (
            .O(N__47099),
            .I(N__47096));
    Span4Mux_v I__10946 (
            .O(N__47096),
            .I(N__47091));
    InMux I__10945 (
            .O(N__47095),
            .I(N__47088));
    InMux I__10944 (
            .O(N__47094),
            .I(N__47085));
    Odrv4 I__10943 (
            .O(N__47091),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__10942 (
            .O(N__47088),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__10941 (
            .O(N__47085),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__10940 (
            .O(N__47078),
            .I(N__47075));
    LocalMux I__10939 (
            .O(N__47075),
            .I(N__47072));
    Odrv12 I__10938 (
            .O(N__47072),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__10937 (
            .O(N__47069),
            .I(N__47063));
    InMux I__10936 (
            .O(N__47068),
            .I(N__47060));
    InMux I__10935 (
            .O(N__47067),
            .I(N__47057));
    InMux I__10934 (
            .O(N__47066),
            .I(N__47054));
    LocalMux I__10933 (
            .O(N__47063),
            .I(N__47051));
    LocalMux I__10932 (
            .O(N__47060),
            .I(N__47048));
    LocalMux I__10931 (
            .O(N__47057),
            .I(N__47045));
    LocalMux I__10930 (
            .O(N__47054),
            .I(N__47042));
    Span12Mux_v I__10929 (
            .O(N__47051),
            .I(N__47037));
    Span12Mux_s10_h I__10928 (
            .O(N__47048),
            .I(N__47037));
    Span4Mux_v I__10927 (
            .O(N__47045),
            .I(N__47034));
    Odrv4 I__10926 (
            .O(N__47042),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv12 I__10925 (
            .O(N__47037),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__10924 (
            .O(N__47034),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__10923 (
            .O(N__47027),
            .I(N__47024));
    LocalMux I__10922 (
            .O(N__47024),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__10921 (
            .O(N__47021),
            .I(N__47018));
    LocalMux I__10920 (
            .O(N__47018),
            .I(N__47015));
    Span4Mux_h I__10919 (
            .O(N__47015),
            .I(N__47012));
    Odrv4 I__10918 (
            .O(N__47012),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    CascadeMux I__10917 (
            .O(N__47009),
            .I(N__47005));
    InMux I__10916 (
            .O(N__47008),
            .I(N__47001));
    InMux I__10915 (
            .O(N__47005),
            .I(N__46996));
    InMux I__10914 (
            .O(N__47004),
            .I(N__46996));
    LocalMux I__10913 (
            .O(N__47001),
            .I(N__46991));
    LocalMux I__10912 (
            .O(N__46996),
            .I(N__46991));
    Span4Mux_h I__10911 (
            .O(N__46991),
            .I(N__46987));
    InMux I__10910 (
            .O(N__46990),
            .I(N__46984));
    Odrv4 I__10909 (
            .O(N__46987),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__10908 (
            .O(N__46984),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__10907 (
            .O(N__46979),
            .I(N__46974));
    InMux I__10906 (
            .O(N__46978),
            .I(N__46969));
    InMux I__10905 (
            .O(N__46977),
            .I(N__46969));
    LocalMux I__10904 (
            .O(N__46974),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__10903 (
            .O(N__46969),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__10902 (
            .O(N__46964),
            .I(N__46956));
    InMux I__10901 (
            .O(N__46963),
            .I(N__46956));
    InMux I__10900 (
            .O(N__46962),
            .I(N__46951));
    InMux I__10899 (
            .O(N__46961),
            .I(N__46951));
    LocalMux I__10898 (
            .O(N__46956),
            .I(N__46948));
    LocalMux I__10897 (
            .O(N__46951),
            .I(N__46945));
    Span4Mux_h I__10896 (
            .O(N__46948),
            .I(N__46942));
    Odrv4 I__10895 (
            .O(N__46945),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__10894 (
            .O(N__46942),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__10893 (
            .O(N__46937),
            .I(N__46934));
    LocalMux I__10892 (
            .O(N__46934),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    CascadeMux I__10891 (
            .O(N__46931),
            .I(N__46927));
    InMux I__10890 (
            .O(N__46930),
            .I(N__46923));
    InMux I__10889 (
            .O(N__46927),
            .I(N__46920));
    InMux I__10888 (
            .O(N__46926),
            .I(N__46917));
    LocalMux I__10887 (
            .O(N__46923),
            .I(N__46914));
    LocalMux I__10886 (
            .O(N__46920),
            .I(N__46911));
    LocalMux I__10885 (
            .O(N__46917),
            .I(N__46908));
    Span4Mux_v I__10884 (
            .O(N__46914),
            .I(N__46905));
    Span4Mux_v I__10883 (
            .O(N__46911),
            .I(N__46901));
    Span4Mux_h I__10882 (
            .O(N__46908),
            .I(N__46896));
    Span4Mux_h I__10881 (
            .O(N__46905),
            .I(N__46896));
    InMux I__10880 (
            .O(N__46904),
            .I(N__46893));
    Odrv4 I__10879 (
            .O(N__46901),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__10878 (
            .O(N__46896),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__10877 (
            .O(N__46893),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__10876 (
            .O(N__46886),
            .I(N__46883));
    LocalMux I__10875 (
            .O(N__46883),
            .I(N__46878));
    InMux I__10874 (
            .O(N__46882),
            .I(N__46875));
    InMux I__10873 (
            .O(N__46881),
            .I(N__46872));
    Odrv4 I__10872 (
            .O(N__46878),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__10871 (
            .O(N__46875),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__10870 (
            .O(N__46872),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__10869 (
            .O(N__46865),
            .I(N__46862));
    LocalMux I__10868 (
            .O(N__46862),
            .I(N__46859));
    Odrv4 I__10867 (
            .O(N__46859),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__10866 (
            .O(N__46856),
            .I(N__46851));
    InMux I__10865 (
            .O(N__46855),
            .I(N__46848));
    InMux I__10864 (
            .O(N__46854),
            .I(N__46845));
    LocalMux I__10863 (
            .O(N__46851),
            .I(N__46842));
    LocalMux I__10862 (
            .O(N__46848),
            .I(N__46839));
    LocalMux I__10861 (
            .O(N__46845),
            .I(N__46836));
    Span4Mux_v I__10860 (
            .O(N__46842),
            .I(N__46833));
    Span4Mux_v I__10859 (
            .O(N__46839),
            .I(N__46829));
    Span4Mux_v I__10858 (
            .O(N__46836),
            .I(N__46824));
    Span4Mux_h I__10857 (
            .O(N__46833),
            .I(N__46824));
    InMux I__10856 (
            .O(N__46832),
            .I(N__46821));
    Odrv4 I__10855 (
            .O(N__46829),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__10854 (
            .O(N__46824),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__10853 (
            .O(N__46821),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__10852 (
            .O(N__46814),
            .I(N__46811));
    LocalMux I__10851 (
            .O(N__46811),
            .I(N__46806));
    InMux I__10850 (
            .O(N__46810),
            .I(N__46803));
    InMux I__10849 (
            .O(N__46809),
            .I(N__46800));
    Odrv12 I__10848 (
            .O(N__46806),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__10847 (
            .O(N__46803),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__10846 (
            .O(N__46800),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__10845 (
            .O(N__46793),
            .I(N__46790));
    LocalMux I__10844 (
            .O(N__46790),
            .I(N__46787));
    Odrv4 I__10843 (
            .O(N__46787),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__10842 (
            .O(N__46784),
            .I(N__46779));
    CascadeMux I__10841 (
            .O(N__46783),
            .I(N__46776));
    InMux I__10840 (
            .O(N__46782),
            .I(N__46773));
    InMux I__10839 (
            .O(N__46779),
            .I(N__46770));
    InMux I__10838 (
            .O(N__46776),
            .I(N__46767));
    LocalMux I__10837 (
            .O(N__46773),
            .I(N__46764));
    LocalMux I__10836 (
            .O(N__46770),
            .I(N__46761));
    LocalMux I__10835 (
            .O(N__46767),
            .I(N__46758));
    Span4Mux_h I__10834 (
            .O(N__46764),
            .I(N__46755));
    Span4Mux_h I__10833 (
            .O(N__46761),
            .I(N__46751));
    Span4Mux_v I__10832 (
            .O(N__46758),
            .I(N__46746));
    Span4Mux_v I__10831 (
            .O(N__46755),
            .I(N__46746));
    InMux I__10830 (
            .O(N__46754),
            .I(N__46743));
    Odrv4 I__10829 (
            .O(N__46751),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10828 (
            .O(N__46746),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__10827 (
            .O(N__46743),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__10826 (
            .O(N__46736),
            .I(N__46733));
    LocalMux I__10825 (
            .O(N__46733),
            .I(N__46728));
    InMux I__10824 (
            .O(N__46732),
            .I(N__46725));
    InMux I__10823 (
            .O(N__46731),
            .I(N__46722));
    Odrv12 I__10822 (
            .O(N__46728),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__10821 (
            .O(N__46725),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__10820 (
            .O(N__46722),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__10819 (
            .O(N__46715),
            .I(N__46712));
    LocalMux I__10818 (
            .O(N__46712),
            .I(N__46709));
    Odrv4 I__10817 (
            .O(N__46709),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__10816 (
            .O(N__46706),
            .I(N__46703));
    InMux I__10815 (
            .O(N__46703),
            .I(N__46698));
    InMux I__10814 (
            .O(N__46702),
            .I(N__46695));
    InMux I__10813 (
            .O(N__46701),
            .I(N__46691));
    LocalMux I__10812 (
            .O(N__46698),
            .I(N__46688));
    LocalMux I__10811 (
            .O(N__46695),
            .I(N__46685));
    InMux I__10810 (
            .O(N__46694),
            .I(N__46682));
    LocalMux I__10809 (
            .O(N__46691),
            .I(N__46679));
    Span4Mux_h I__10808 (
            .O(N__46688),
            .I(N__46676));
    Span4Mux_v I__10807 (
            .O(N__46685),
            .I(N__46673));
    LocalMux I__10806 (
            .O(N__46682),
            .I(N__46670));
    Span4Mux_h I__10805 (
            .O(N__46679),
            .I(N__46667));
    Span4Mux_v I__10804 (
            .O(N__46676),
            .I(N__46664));
    Span4Mux_h I__10803 (
            .O(N__46673),
            .I(N__46661));
    Span12Mux_v I__10802 (
            .O(N__46670),
            .I(N__46658));
    Odrv4 I__10801 (
            .O(N__46667),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10800 (
            .O(N__46664),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10799 (
            .O(N__46661),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv12 I__10798 (
            .O(N__46658),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__10797 (
            .O(N__46649),
            .I(N__46645));
    CascadeMux I__10796 (
            .O(N__46648),
            .I(N__46642));
    LocalMux I__10795 (
            .O(N__46645),
            .I(N__46639));
    InMux I__10794 (
            .O(N__46642),
            .I(N__46635));
    Span4Mux_h I__10793 (
            .O(N__46639),
            .I(N__46632));
    InMux I__10792 (
            .O(N__46638),
            .I(N__46629));
    LocalMux I__10791 (
            .O(N__46635),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__10790 (
            .O(N__46632),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__10789 (
            .O(N__46629),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__10788 (
            .O(N__46622),
            .I(N__46619));
    LocalMux I__10787 (
            .O(N__46619),
            .I(N__46616));
    Odrv12 I__10786 (
            .O(N__46616),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__10785 (
            .O(N__46613),
            .I(N__46606));
    InMux I__10784 (
            .O(N__46612),
            .I(N__46606));
    InMux I__10783 (
            .O(N__46611),
            .I(N__46603));
    LocalMux I__10782 (
            .O(N__46606),
            .I(N__46600));
    LocalMux I__10781 (
            .O(N__46603),
            .I(N__46597));
    Span4Mux_h I__10780 (
            .O(N__46600),
            .I(N__46594));
    Span4Mux_h I__10779 (
            .O(N__46597),
            .I(N__46588));
    Span4Mux_v I__10778 (
            .O(N__46594),
            .I(N__46588));
    InMux I__10777 (
            .O(N__46593),
            .I(N__46585));
    Odrv4 I__10776 (
            .O(N__46588),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__10775 (
            .O(N__46585),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__10774 (
            .O(N__46580),
            .I(N__46573));
    InMux I__10773 (
            .O(N__46579),
            .I(N__46573));
    InMux I__10772 (
            .O(N__46578),
            .I(N__46570));
    LocalMux I__10771 (
            .O(N__46573),
            .I(N__46567));
    LocalMux I__10770 (
            .O(N__46570),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__10769 (
            .O(N__46567),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__10768 (
            .O(N__46562),
            .I(N__46559));
    LocalMux I__10767 (
            .O(N__46559),
            .I(N__46556));
    Span4Mux_h I__10766 (
            .O(N__46556),
            .I(N__46553));
    Odrv4 I__10765 (
            .O(N__46553),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    CascadeMux I__10764 (
            .O(N__46550),
            .I(N__46547));
    InMux I__10763 (
            .O(N__46547),
            .I(N__46542));
    InMux I__10762 (
            .O(N__46546),
            .I(N__46539));
    InMux I__10761 (
            .O(N__46545),
            .I(N__46536));
    LocalMux I__10760 (
            .O(N__46542),
            .I(N__46533));
    LocalMux I__10759 (
            .O(N__46539),
            .I(N__46530));
    LocalMux I__10758 (
            .O(N__46536),
            .I(N__46527));
    Span4Mux_v I__10757 (
            .O(N__46533),
            .I(N__46522));
    Span4Mux_h I__10756 (
            .O(N__46530),
            .I(N__46522));
    Span4Mux_v I__10755 (
            .O(N__46527),
            .I(N__46518));
    Span4Mux_v I__10754 (
            .O(N__46522),
            .I(N__46515));
    InMux I__10753 (
            .O(N__46521),
            .I(N__46512));
    Odrv4 I__10752 (
            .O(N__46518),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__10751 (
            .O(N__46515),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__10750 (
            .O(N__46512),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__10749 (
            .O(N__46505),
            .I(N__46502));
    LocalMux I__10748 (
            .O(N__46502),
            .I(N__46497));
    InMux I__10747 (
            .O(N__46501),
            .I(N__46494));
    InMux I__10746 (
            .O(N__46500),
            .I(N__46491));
    Odrv4 I__10745 (
            .O(N__46497),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__10744 (
            .O(N__46494),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__10743 (
            .O(N__46491),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__10742 (
            .O(N__46484),
            .I(N__46481));
    LocalMux I__10741 (
            .O(N__46481),
            .I(N__46478));
    Odrv4 I__10740 (
            .O(N__46478),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__10739 (
            .O(N__46475),
            .I(N__46472));
    LocalMux I__10738 (
            .O(N__46472),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__10737 (
            .O(N__46469),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__10736 (
            .O(N__46466),
            .I(N__46463));
    InMux I__10735 (
            .O(N__46463),
            .I(N__46456));
    InMux I__10734 (
            .O(N__46462),
            .I(N__46453));
    InMux I__10733 (
            .O(N__46461),
            .I(N__46446));
    InMux I__10732 (
            .O(N__46460),
            .I(N__46446));
    InMux I__10731 (
            .O(N__46459),
            .I(N__46446));
    LocalMux I__10730 (
            .O(N__46456),
            .I(N__46433));
    LocalMux I__10729 (
            .O(N__46453),
            .I(N__46433));
    LocalMux I__10728 (
            .O(N__46446),
            .I(N__46430));
    InMux I__10727 (
            .O(N__46445),
            .I(N__46413));
    InMux I__10726 (
            .O(N__46444),
            .I(N__46413));
    InMux I__10725 (
            .O(N__46443),
            .I(N__46413));
    InMux I__10724 (
            .O(N__46442),
            .I(N__46413));
    InMux I__10723 (
            .O(N__46441),
            .I(N__46413));
    InMux I__10722 (
            .O(N__46440),
            .I(N__46413));
    InMux I__10721 (
            .O(N__46439),
            .I(N__46413));
    InMux I__10720 (
            .O(N__46438),
            .I(N__46413));
    Span4Mux_v I__10719 (
            .O(N__46433),
            .I(N__46406));
    Span4Mux_v I__10718 (
            .O(N__46430),
            .I(N__46406));
    LocalMux I__10717 (
            .O(N__46413),
            .I(N__46406));
    Odrv4 I__10716 (
            .O(N__46406),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__10715 (
            .O(N__46403),
            .I(N__46400));
    LocalMux I__10714 (
            .O(N__46400),
            .I(N__46397));
    Odrv12 I__10713 (
            .O(N__46397),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__10712 (
            .O(N__46394),
            .I(N__46390));
    CascadeMux I__10711 (
            .O(N__46393),
            .I(N__46387));
    LocalMux I__10710 (
            .O(N__46390),
            .I(N__46384));
    InMux I__10709 (
            .O(N__46387),
            .I(N__46381));
    Span4Mux_h I__10708 (
            .O(N__46384),
            .I(N__46377));
    LocalMux I__10707 (
            .O(N__46381),
            .I(N__46374));
    InMux I__10706 (
            .O(N__46380),
            .I(N__46371));
    Span4Mux_v I__10705 (
            .O(N__46377),
            .I(N__46366));
    Span4Mux_h I__10704 (
            .O(N__46374),
            .I(N__46366));
    LocalMux I__10703 (
            .O(N__46371),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__10702 (
            .O(N__46366),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__10701 (
            .O(N__46361),
            .I(N__46358));
    LocalMux I__10700 (
            .O(N__46358),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__10699 (
            .O(N__46355),
            .I(N__46350));
    CascadeMux I__10698 (
            .O(N__46354),
            .I(N__46346));
    InMux I__10697 (
            .O(N__46353),
            .I(N__46341));
    InMux I__10696 (
            .O(N__46350),
            .I(N__46341));
    CascadeMux I__10695 (
            .O(N__46349),
            .I(N__46338));
    InMux I__10694 (
            .O(N__46346),
            .I(N__46335));
    LocalMux I__10693 (
            .O(N__46341),
            .I(N__46332));
    InMux I__10692 (
            .O(N__46338),
            .I(N__46329));
    LocalMux I__10691 (
            .O(N__46335),
            .I(N__46326));
    Odrv12 I__10690 (
            .O(N__46332),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__10689 (
            .O(N__46329),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__10688 (
            .O(N__46326),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__10687 (
            .O(N__46319),
            .I(N__46316));
    LocalMux I__10686 (
            .O(N__46316),
            .I(N__46313));
    Span4Mux_h I__10685 (
            .O(N__46313),
            .I(N__46310));
    Odrv4 I__10684 (
            .O(N__46310),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__10683 (
            .O(N__46307),
            .I(N__46304));
    InMux I__10682 (
            .O(N__46304),
            .I(N__46295));
    InMux I__10681 (
            .O(N__46303),
            .I(N__46295));
    InMux I__10680 (
            .O(N__46302),
            .I(N__46295));
    LocalMux I__10679 (
            .O(N__46295),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__10678 (
            .O(N__46292),
            .I(N__46280));
    InMux I__10677 (
            .O(N__46291),
            .I(N__46280));
    InMux I__10676 (
            .O(N__46290),
            .I(N__46280));
    InMux I__10675 (
            .O(N__46289),
            .I(N__46280));
    LocalMux I__10674 (
            .O(N__46280),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__10673 (
            .O(N__46277),
            .I(N__46274));
    LocalMux I__10672 (
            .O(N__46274),
            .I(N__46271));
    Odrv12 I__10671 (
            .O(N__46271),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    CascadeMux I__10670 (
            .O(N__46268),
            .I(N__46263));
    CascadeMux I__10669 (
            .O(N__46267),
            .I(N__46260));
    InMux I__10668 (
            .O(N__46266),
            .I(N__46257));
    InMux I__10667 (
            .O(N__46263),
            .I(N__46254));
    InMux I__10666 (
            .O(N__46260),
            .I(N__46251));
    LocalMux I__10665 (
            .O(N__46257),
            .I(N__46248));
    LocalMux I__10664 (
            .O(N__46254),
            .I(N__46245));
    LocalMux I__10663 (
            .O(N__46251),
            .I(N__46242));
    Span4Mux_h I__10662 (
            .O(N__46248),
            .I(N__46239));
    Span4Mux_v I__10661 (
            .O(N__46245),
            .I(N__46233));
    Span4Mux_v I__10660 (
            .O(N__46242),
            .I(N__46233));
    Span4Mux_v I__10659 (
            .O(N__46239),
            .I(N__46230));
    InMux I__10658 (
            .O(N__46238),
            .I(N__46227));
    Odrv4 I__10657 (
            .O(N__46233),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__10656 (
            .O(N__46230),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__10655 (
            .O(N__46227),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__10654 (
            .O(N__46220),
            .I(N__46215));
    InMux I__10653 (
            .O(N__46219),
            .I(N__46212));
    InMux I__10652 (
            .O(N__46218),
            .I(N__46209));
    LocalMux I__10651 (
            .O(N__46215),
            .I(N__46206));
    LocalMux I__10650 (
            .O(N__46212),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__10649 (
            .O(N__46209),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__10648 (
            .O(N__46206),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__10647 (
            .O(N__46199),
            .I(N__46196));
    LocalMux I__10646 (
            .O(N__46196),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__10645 (
            .O(N__46193),
            .I(N__46187));
    InMux I__10644 (
            .O(N__46192),
            .I(N__46187));
    LocalMux I__10643 (
            .O(N__46187),
            .I(N__46184));
    Span4Mux_h I__10642 (
            .O(N__46184),
            .I(N__46180));
    InMux I__10641 (
            .O(N__46183),
            .I(N__46177));
    Odrv4 I__10640 (
            .O(N__46180),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__10639 (
            .O(N__46177),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__10638 (
            .O(N__46172),
            .I(N__46169));
    LocalMux I__10637 (
            .O(N__46169),
            .I(N__46166));
    Span4Mux_v I__10636 (
            .O(N__46166),
            .I(N__46163));
    Odrv4 I__10635 (
            .O(N__46163),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__10634 (
            .O(N__46160),
            .I(N__46157));
    InMux I__10633 (
            .O(N__46157),
            .I(N__46154));
    LocalMux I__10632 (
            .O(N__46154),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__10631 (
            .O(N__46151),
            .I(N__46142));
    CascadeMux I__10630 (
            .O(N__46150),
            .I(N__46139));
    CascadeMux I__10629 (
            .O(N__46149),
            .I(N__46136));
    CascadeMux I__10628 (
            .O(N__46148),
            .I(N__46133));
    CascadeMux I__10627 (
            .O(N__46147),
            .I(N__46130));
    CascadeMux I__10626 (
            .O(N__46146),
            .I(N__46126));
    CascadeMux I__10625 (
            .O(N__46145),
            .I(N__46123));
    InMux I__10624 (
            .O(N__46142),
            .I(N__46104));
    InMux I__10623 (
            .O(N__46139),
            .I(N__46104));
    InMux I__10622 (
            .O(N__46136),
            .I(N__46104));
    InMux I__10621 (
            .O(N__46133),
            .I(N__46104));
    InMux I__10620 (
            .O(N__46130),
            .I(N__46095));
    InMux I__10619 (
            .O(N__46129),
            .I(N__46095));
    InMux I__10618 (
            .O(N__46126),
            .I(N__46095));
    InMux I__10617 (
            .O(N__46123),
            .I(N__46095));
    CascadeMux I__10616 (
            .O(N__46122),
            .I(N__46091));
    CascadeMux I__10615 (
            .O(N__46121),
            .I(N__46088));
    CascadeMux I__10614 (
            .O(N__46120),
            .I(N__46085));
    CascadeMux I__10613 (
            .O(N__46119),
            .I(N__46082));
    CascadeMux I__10612 (
            .O(N__46118),
            .I(N__46078));
    CascadeMux I__10611 (
            .O(N__46117),
            .I(N__46075));
    CascadeMux I__10610 (
            .O(N__46116),
            .I(N__46072));
    CascadeMux I__10609 (
            .O(N__46115),
            .I(N__46069));
    CascadeMux I__10608 (
            .O(N__46114),
            .I(N__46065));
    CascadeMux I__10607 (
            .O(N__46113),
            .I(N__46062));
    LocalMux I__10606 (
            .O(N__46104),
            .I(N__46056));
    LocalMux I__10605 (
            .O(N__46095),
            .I(N__46053));
    InMux I__10604 (
            .O(N__46094),
            .I(N__46042));
    InMux I__10603 (
            .O(N__46091),
            .I(N__46042));
    InMux I__10602 (
            .O(N__46088),
            .I(N__46042));
    InMux I__10601 (
            .O(N__46085),
            .I(N__46042));
    InMux I__10600 (
            .O(N__46082),
            .I(N__46042));
    InMux I__10599 (
            .O(N__46081),
            .I(N__46032));
    InMux I__10598 (
            .O(N__46078),
            .I(N__46017));
    InMux I__10597 (
            .O(N__46075),
            .I(N__46017));
    InMux I__10596 (
            .O(N__46072),
            .I(N__46017));
    InMux I__10595 (
            .O(N__46069),
            .I(N__46008));
    InMux I__10594 (
            .O(N__46068),
            .I(N__46008));
    InMux I__10593 (
            .O(N__46065),
            .I(N__46008));
    InMux I__10592 (
            .O(N__46062),
            .I(N__46008));
    CascadeMux I__10591 (
            .O(N__46061),
            .I(N__46005));
    CascadeMux I__10590 (
            .O(N__46060),
            .I(N__46002));
    CascadeMux I__10589 (
            .O(N__46059),
            .I(N__45999));
    Span4Mux_v I__10588 (
            .O(N__46056),
            .I(N__45992));
    Span4Mux_h I__10587 (
            .O(N__46053),
            .I(N__45992));
    LocalMux I__10586 (
            .O(N__46042),
            .I(N__45992));
    CascadeMux I__10585 (
            .O(N__46041),
            .I(N__45989));
    CascadeMux I__10584 (
            .O(N__46040),
            .I(N__45986));
    CascadeMux I__10583 (
            .O(N__46039),
            .I(N__45983));
    CascadeMux I__10582 (
            .O(N__46038),
            .I(N__45980));
    CascadeMux I__10581 (
            .O(N__46037),
            .I(N__45977));
    CascadeMux I__10580 (
            .O(N__46036),
            .I(N__45974));
    CascadeMux I__10579 (
            .O(N__46035),
            .I(N__45971));
    LocalMux I__10578 (
            .O(N__46032),
            .I(N__45968));
    InMux I__10577 (
            .O(N__46031),
            .I(N__45963));
    InMux I__10576 (
            .O(N__46030),
            .I(N__45956));
    InMux I__10575 (
            .O(N__46029),
            .I(N__45956));
    InMux I__10574 (
            .O(N__46028),
            .I(N__45956));
    InMux I__10573 (
            .O(N__46027),
            .I(N__45947));
    InMux I__10572 (
            .O(N__46026),
            .I(N__45947));
    InMux I__10571 (
            .O(N__46025),
            .I(N__45947));
    InMux I__10570 (
            .O(N__46024),
            .I(N__45947));
    LocalMux I__10569 (
            .O(N__46017),
            .I(N__45942));
    LocalMux I__10568 (
            .O(N__46008),
            .I(N__45942));
    InMux I__10567 (
            .O(N__46005),
            .I(N__45935));
    InMux I__10566 (
            .O(N__46002),
            .I(N__45935));
    InMux I__10565 (
            .O(N__45999),
            .I(N__45935));
    Span4Mux_v I__10564 (
            .O(N__45992),
            .I(N__45932));
    InMux I__10563 (
            .O(N__45989),
            .I(N__45925));
    InMux I__10562 (
            .O(N__45986),
            .I(N__45925));
    InMux I__10561 (
            .O(N__45983),
            .I(N__45925));
    InMux I__10560 (
            .O(N__45980),
            .I(N__45916));
    InMux I__10559 (
            .O(N__45977),
            .I(N__45916));
    InMux I__10558 (
            .O(N__45974),
            .I(N__45916));
    InMux I__10557 (
            .O(N__45971),
            .I(N__45916));
    Span4Mux_v I__10556 (
            .O(N__45968),
            .I(N__45913));
    InMux I__10555 (
            .O(N__45967),
            .I(N__45909));
    CascadeMux I__10554 (
            .O(N__45966),
            .I(N__45904));
    LocalMux I__10553 (
            .O(N__45963),
            .I(N__45897));
    LocalMux I__10552 (
            .O(N__45956),
            .I(N__45897));
    LocalMux I__10551 (
            .O(N__45947),
            .I(N__45897));
    Span4Mux_v I__10550 (
            .O(N__45942),
            .I(N__45878));
    LocalMux I__10549 (
            .O(N__45935),
            .I(N__45878));
    Span4Mux_v I__10548 (
            .O(N__45932),
            .I(N__45878));
    LocalMux I__10547 (
            .O(N__45925),
            .I(N__45878));
    LocalMux I__10546 (
            .O(N__45916),
            .I(N__45878));
    Span4Mux_h I__10545 (
            .O(N__45913),
            .I(N__45875));
    InMux I__10544 (
            .O(N__45912),
            .I(N__45872));
    LocalMux I__10543 (
            .O(N__45909),
            .I(N__45869));
    InMux I__10542 (
            .O(N__45908),
            .I(N__45866));
    InMux I__10541 (
            .O(N__45907),
            .I(N__45861));
    InMux I__10540 (
            .O(N__45904),
            .I(N__45861));
    Span4Mux_v I__10539 (
            .O(N__45897),
            .I(N__45858));
    InMux I__10538 (
            .O(N__45896),
            .I(N__45849));
    InMux I__10537 (
            .O(N__45895),
            .I(N__45849));
    InMux I__10536 (
            .O(N__45894),
            .I(N__45849));
    InMux I__10535 (
            .O(N__45893),
            .I(N__45840));
    InMux I__10534 (
            .O(N__45892),
            .I(N__45840));
    InMux I__10533 (
            .O(N__45891),
            .I(N__45840));
    InMux I__10532 (
            .O(N__45890),
            .I(N__45840));
    CascadeMux I__10531 (
            .O(N__45889),
            .I(N__45837));
    Sp12to4 I__10530 (
            .O(N__45878),
            .I(N__45833));
    Span4Mux_v I__10529 (
            .O(N__45875),
            .I(N__45830));
    LocalMux I__10528 (
            .O(N__45872),
            .I(N__45825));
    Span4Mux_s1_v I__10527 (
            .O(N__45869),
            .I(N__45825));
    LocalMux I__10526 (
            .O(N__45866),
            .I(N__45822));
    LocalMux I__10525 (
            .O(N__45861),
            .I(N__45819));
    Span4Mux_v I__10524 (
            .O(N__45858),
            .I(N__45816));
    InMux I__10523 (
            .O(N__45857),
            .I(N__45813));
    CascadeMux I__10522 (
            .O(N__45856),
            .I(N__45810));
    LocalMux I__10521 (
            .O(N__45849),
            .I(N__45805));
    LocalMux I__10520 (
            .O(N__45840),
            .I(N__45805));
    InMux I__10519 (
            .O(N__45837),
            .I(N__45800));
    InMux I__10518 (
            .O(N__45836),
            .I(N__45800));
    Span12Mux_v I__10517 (
            .O(N__45833),
            .I(N__45795));
    Sp12to4 I__10516 (
            .O(N__45830),
            .I(N__45795));
    Span4Mux_v I__10515 (
            .O(N__45825),
            .I(N__45790));
    Span4Mux_v I__10514 (
            .O(N__45822),
            .I(N__45790));
    Span12Mux_v I__10513 (
            .O(N__45819),
            .I(N__45787));
    Sp12to4 I__10512 (
            .O(N__45816),
            .I(N__45782));
    LocalMux I__10511 (
            .O(N__45813),
            .I(N__45782));
    InMux I__10510 (
            .O(N__45810),
            .I(N__45779));
    Span4Mux_s2_h I__10509 (
            .O(N__45805),
            .I(N__45774));
    LocalMux I__10508 (
            .O(N__45800),
            .I(N__45774));
    Span12Mux_h I__10507 (
            .O(N__45795),
            .I(N__45771));
    Span4Mux_v I__10506 (
            .O(N__45790),
            .I(N__45768));
    Span12Mux_h I__10505 (
            .O(N__45787),
            .I(N__45759));
    Span12Mux_s2_h I__10504 (
            .O(N__45782),
            .I(N__45759));
    LocalMux I__10503 (
            .O(N__45779),
            .I(N__45759));
    Sp12to4 I__10502 (
            .O(N__45774),
            .I(N__45759));
    Odrv12 I__10501 (
            .O(N__45771),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10500 (
            .O(N__45768),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10499 (
            .O(N__45759),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__10498 (
            .O(N__45752),
            .I(N__45749));
    InMux I__10497 (
            .O(N__45749),
            .I(N__45746));
    LocalMux I__10496 (
            .O(N__45746),
            .I(N__45743));
    Odrv4 I__10495 (
            .O(N__45743),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__10494 (
            .O(N__45740),
            .I(N__45737));
    LocalMux I__10493 (
            .O(N__45737),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__10492 (
            .O(N__45734),
            .I(N__45731));
    LocalMux I__10491 (
            .O(N__45731),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__10490 (
            .O(N__45728),
            .I(N__45725));
    LocalMux I__10489 (
            .O(N__45725),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__10488 (
            .O(N__45722),
            .I(N__45719));
    LocalMux I__10487 (
            .O(N__45719),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__10486 (
            .O(N__45716),
            .I(N__45713));
    LocalMux I__10485 (
            .O(N__45713),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__10484 (
            .O(N__45710),
            .I(N__45707));
    LocalMux I__10483 (
            .O(N__45707),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__10482 (
            .O(N__45704),
            .I(N__45701));
    InMux I__10481 (
            .O(N__45701),
            .I(N__45698));
    LocalMux I__10480 (
            .O(N__45698),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__10479 (
            .O(N__45695),
            .I(N__45692));
    LocalMux I__10478 (
            .O(N__45692),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__10477 (
            .O(N__45689),
            .I(N__45686));
    LocalMux I__10476 (
            .O(N__45686),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__10475 (
            .O(N__45683),
            .I(N__45680));
    LocalMux I__10474 (
            .O(N__45680),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__10473 (
            .O(N__45677),
            .I(N__45674));
    LocalMux I__10472 (
            .O(N__45674),
            .I(N__45671));
    Odrv12 I__10471 (
            .O(N__45671),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__10470 (
            .O(N__45668),
            .I(N__45663));
    InMux I__10469 (
            .O(N__45667),
            .I(N__45660));
    InMux I__10468 (
            .O(N__45666),
            .I(N__45657));
    LocalMux I__10467 (
            .O(N__45663),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__10466 (
            .O(N__45660),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__10465 (
            .O(N__45657),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__10464 (
            .O(N__45650),
            .I(N__45646));
    InMux I__10463 (
            .O(N__45649),
            .I(N__45643));
    InMux I__10462 (
            .O(N__45646),
            .I(N__45640));
    LocalMux I__10461 (
            .O(N__45643),
            .I(N__45637));
    LocalMux I__10460 (
            .O(N__45640),
            .I(N__45634));
    Span4Mux_h I__10459 (
            .O(N__45637),
            .I(N__45631));
    Span4Mux_v I__10458 (
            .O(N__45634),
            .I(N__45628));
    Span4Mux_h I__10457 (
            .O(N__45631),
            .I(N__45625));
    Span4Mux_h I__10456 (
            .O(N__45628),
            .I(N__45622));
    Odrv4 I__10455 (
            .O(N__45625),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    Odrv4 I__10454 (
            .O(N__45622),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    InMux I__10453 (
            .O(N__45617),
            .I(N__45612));
    InMux I__10452 (
            .O(N__45616),
            .I(N__45609));
    InMux I__10451 (
            .O(N__45615),
            .I(N__45606));
    LocalMux I__10450 (
            .O(N__45612),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10449 (
            .O(N__45609),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10448 (
            .O(N__45606),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__10447 (
            .O(N__45599),
            .I(N__45596));
    LocalMux I__10446 (
            .O(N__45596),
            .I(N__45591));
    InMux I__10445 (
            .O(N__45595),
            .I(N__45588));
    InMux I__10444 (
            .O(N__45594),
            .I(N__45585));
    Span4Mux_h I__10443 (
            .O(N__45591),
            .I(N__45580));
    LocalMux I__10442 (
            .O(N__45588),
            .I(N__45580));
    LocalMux I__10441 (
            .O(N__45585),
            .I(N__45577));
    Span4Mux_h I__10440 (
            .O(N__45580),
            .I(N__45574));
    Odrv12 I__10439 (
            .O(N__45577),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__10438 (
            .O(N__45574),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    CEMux I__10437 (
            .O(N__45569),
            .I(N__45551));
    CEMux I__10436 (
            .O(N__45568),
            .I(N__45551));
    CEMux I__10435 (
            .O(N__45567),
            .I(N__45551));
    CEMux I__10434 (
            .O(N__45566),
            .I(N__45551));
    CEMux I__10433 (
            .O(N__45565),
            .I(N__45551));
    CEMux I__10432 (
            .O(N__45564),
            .I(N__45551));
    GlobalMux I__10431 (
            .O(N__45551),
            .I(N__45548));
    gio2CtrlBuf I__10430 (
            .O(N__45548),
            .I(\delay_measurement_inst.delay_tr_timer.N_304_i_g ));
    InMux I__10429 (
            .O(N__45545),
            .I(N__45542));
    LocalMux I__10428 (
            .O(N__45542),
            .I(N__45538));
    InMux I__10427 (
            .O(N__45541),
            .I(N__45535));
    Span4Mux_s1_v I__10426 (
            .O(N__45538),
            .I(N__45530));
    LocalMux I__10425 (
            .O(N__45535),
            .I(N__45530));
    Span4Mux_v I__10424 (
            .O(N__45530),
            .I(N__45527));
    Span4Mux_h I__10423 (
            .O(N__45527),
            .I(N__45524));
    Sp12to4 I__10422 (
            .O(N__45524),
            .I(N__45520));
    InMux I__10421 (
            .O(N__45523),
            .I(N__45517));
    Span12Mux_v I__10420 (
            .O(N__45520),
            .I(N__45514));
    LocalMux I__10419 (
            .O(N__45517),
            .I(N__45511));
    Span12Mux_v I__10418 (
            .O(N__45514),
            .I(N__45507));
    Span12Mux_h I__10417 (
            .O(N__45511),
            .I(N__45504));
    InMux I__10416 (
            .O(N__45510),
            .I(N__45501));
    Span12Mux_h I__10415 (
            .O(N__45507),
            .I(N__45496));
    Span12Mux_v I__10414 (
            .O(N__45504),
            .I(N__45496));
    LocalMux I__10413 (
            .O(N__45501),
            .I(N__45493));
    Odrv12 I__10412 (
            .O(N__45496),
            .I(start_stop_c));
    Odrv12 I__10411 (
            .O(N__45493),
            .I(start_stop_c));
    InMux I__10410 (
            .O(N__45488),
            .I(N__45483));
    InMux I__10409 (
            .O(N__45487),
            .I(N__45476));
    InMux I__10408 (
            .O(N__45486),
            .I(N__45476));
    LocalMux I__10407 (
            .O(N__45483),
            .I(N__45473));
    InMux I__10406 (
            .O(N__45482),
            .I(N__45470));
    InMux I__10405 (
            .O(N__45481),
            .I(N__45467));
    LocalMux I__10404 (
            .O(N__45476),
            .I(N__45464));
    Span4Mux_v I__10403 (
            .O(N__45473),
            .I(N__45459));
    LocalMux I__10402 (
            .O(N__45470),
            .I(N__45459));
    LocalMux I__10401 (
            .O(N__45467),
            .I(N__45455));
    Span4Mux_h I__10400 (
            .O(N__45464),
            .I(N__45452));
    Span4Mux_v I__10399 (
            .O(N__45459),
            .I(N__45449));
    InMux I__10398 (
            .O(N__45458),
            .I(N__45446));
    Span4Mux_v I__10397 (
            .O(N__45455),
            .I(N__45439));
    Span4Mux_v I__10396 (
            .O(N__45452),
            .I(N__45439));
    Span4Mux_h I__10395 (
            .O(N__45449),
            .I(N__45439));
    LocalMux I__10394 (
            .O(N__45446),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__10393 (
            .O(N__45439),
            .I(phase_controller_inst1_state_4));
    InMux I__10392 (
            .O(N__45434),
            .I(N__45430));
    InMux I__10391 (
            .O(N__45433),
            .I(N__45427));
    LocalMux I__10390 (
            .O(N__45430),
            .I(N__45424));
    LocalMux I__10389 (
            .O(N__45427),
            .I(N__45421));
    Span4Mux_v I__10388 (
            .O(N__45424),
            .I(N__45418));
    Span4Mux_h I__10387 (
            .O(N__45421),
            .I(N__45415));
    Span4Mux_v I__10386 (
            .O(N__45418),
            .I(N__45412));
    Span4Mux_v I__10385 (
            .O(N__45415),
            .I(N__45409));
    Odrv4 I__10384 (
            .O(N__45412),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__10383 (
            .O(N__45409),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    CascadeMux I__10382 (
            .O(N__45404),
            .I(N__45401));
    InMux I__10381 (
            .O(N__45401),
            .I(N__45398));
    LocalMux I__10380 (
            .O(N__45398),
            .I(N__45393));
    InMux I__10379 (
            .O(N__45397),
            .I(N__45388));
    InMux I__10378 (
            .O(N__45396),
            .I(N__45388));
    Span4Mux_v I__10377 (
            .O(N__45393),
            .I(N__45385));
    LocalMux I__10376 (
            .O(N__45388),
            .I(N__45382));
    Odrv4 I__10375 (
            .O(N__45385),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__10374 (
            .O(N__45382),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__10373 (
            .O(N__45377),
            .I(N__45374));
    LocalMux I__10372 (
            .O(N__45374),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__10371 (
            .O(N__45371),
            .I(N__45368));
    LocalMux I__10370 (
            .O(N__45368),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__10369 (
            .O(N__45365),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__10368 (
            .O(N__45362),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__10367 (
            .O(N__45359),
            .I(N__45356));
    InMux I__10366 (
            .O(N__45356),
            .I(N__45353));
    LocalMux I__10365 (
            .O(N__45353),
            .I(N__45350));
    Span4Mux_h I__10364 (
            .O(N__45350),
            .I(N__45347));
    Span4Mux_v I__10363 (
            .O(N__45347),
            .I(N__45344));
    Odrv4 I__10362 (
            .O(N__45344),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__10361 (
            .O(N__45341),
            .I(N__45338));
    InMux I__10360 (
            .O(N__45338),
            .I(N__45335));
    LocalMux I__10359 (
            .O(N__45335),
            .I(N__45332));
    Span4Mux_h I__10358 (
            .O(N__45332),
            .I(N__45329));
    Odrv4 I__10357 (
            .O(N__45329),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    CascadeMux I__10356 (
            .O(N__45326),
            .I(N__45321));
    InMux I__10355 (
            .O(N__45325),
            .I(N__45318));
    InMux I__10354 (
            .O(N__45324),
            .I(N__45315));
    InMux I__10353 (
            .O(N__45321),
            .I(N__45312));
    LocalMux I__10352 (
            .O(N__45318),
            .I(N__45309));
    LocalMux I__10351 (
            .O(N__45315),
            .I(N__45306));
    LocalMux I__10350 (
            .O(N__45312),
            .I(N__45303));
    Span4Mux_h I__10349 (
            .O(N__45309),
            .I(N__45300));
    Span4Mux_h I__10348 (
            .O(N__45306),
            .I(N__45295));
    Span4Mux_h I__10347 (
            .O(N__45303),
            .I(N__45295));
    Odrv4 I__10346 (
            .O(N__45300),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__10345 (
            .O(N__45295),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__10344 (
            .O(N__45290),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    CascadeMux I__10343 (
            .O(N__45287),
            .I(N__45284));
    InMux I__10342 (
            .O(N__45284),
            .I(N__45278));
    InMux I__10341 (
            .O(N__45283),
            .I(N__45273));
    InMux I__10340 (
            .O(N__45282),
            .I(N__45273));
    InMux I__10339 (
            .O(N__45281),
            .I(N__45270));
    LocalMux I__10338 (
            .O(N__45278),
            .I(N__45267));
    LocalMux I__10337 (
            .O(N__45273),
            .I(N__45264));
    LocalMux I__10336 (
            .O(N__45270),
            .I(N__45261));
    Span4Mux_v I__10335 (
            .O(N__45267),
            .I(N__45258));
    Span12Mux_s10_h I__10334 (
            .O(N__45264),
            .I(N__45255));
    Span4Mux_h I__10333 (
            .O(N__45261),
            .I(N__45252));
    Odrv4 I__10332 (
            .O(N__45258),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv12 I__10331 (
            .O(N__45255),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10330 (
            .O(N__45252),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10329 (
            .O(N__45245),
            .I(N__45242));
    LocalMux I__10328 (
            .O(N__45242),
            .I(N__45239));
    Odrv4 I__10327 (
            .O(N__45239),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__10326 (
            .O(N__45236),
            .I(N__45233));
    LocalMux I__10325 (
            .O(N__45233),
            .I(N__45228));
    InMux I__10324 (
            .O(N__45232),
            .I(N__45222));
    InMux I__10323 (
            .O(N__45231),
            .I(N__45222));
    Span4Mux_v I__10322 (
            .O(N__45228),
            .I(N__45219));
    InMux I__10321 (
            .O(N__45227),
            .I(N__45216));
    LocalMux I__10320 (
            .O(N__45222),
            .I(N__45213));
    Span4Mux_v I__10319 (
            .O(N__45219),
            .I(N__45210));
    LocalMux I__10318 (
            .O(N__45216),
            .I(N__45207));
    Odrv12 I__10317 (
            .O(N__45213),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__10316 (
            .O(N__45210),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__10315 (
            .O(N__45207),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__10314 (
            .O(N__45200),
            .I(N__45197));
    LocalMux I__10313 (
            .O(N__45197),
            .I(N__45194));
    Odrv12 I__10312 (
            .O(N__45194),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    CascadeMux I__10311 (
            .O(N__45191),
            .I(N__45186));
    InMux I__10310 (
            .O(N__45190),
            .I(N__45183));
    InMux I__10309 (
            .O(N__45189),
            .I(N__45180));
    InMux I__10308 (
            .O(N__45186),
            .I(N__45177));
    LocalMux I__10307 (
            .O(N__45183),
            .I(N__45172));
    LocalMux I__10306 (
            .O(N__45180),
            .I(N__45172));
    LocalMux I__10305 (
            .O(N__45177),
            .I(N__45168));
    Span4Mux_v I__10304 (
            .O(N__45172),
            .I(N__45165));
    InMux I__10303 (
            .O(N__45171),
            .I(N__45162));
    Span4Mux_h I__10302 (
            .O(N__45168),
            .I(N__45159));
    Span4Mux_v I__10301 (
            .O(N__45165),
            .I(N__45154));
    LocalMux I__10300 (
            .O(N__45162),
            .I(N__45154));
    Odrv4 I__10299 (
            .O(N__45159),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__10298 (
            .O(N__45154),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__10297 (
            .O(N__45149),
            .I(N__45146));
    LocalMux I__10296 (
            .O(N__45146),
            .I(N__45143));
    Odrv12 I__10295 (
            .O(N__45143),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__10294 (
            .O(N__45140),
            .I(N__45137));
    LocalMux I__10293 (
            .O(N__45137),
            .I(N__45134));
    Odrv4 I__10292 (
            .O(N__45134),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__10291 (
            .O(N__45131),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__10290 (
            .O(N__45128),
            .I(N__45125));
    LocalMux I__10289 (
            .O(N__45125),
            .I(N__45122));
    Odrv4 I__10288 (
            .O(N__45122),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__10287 (
            .O(N__45119),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__10286 (
            .O(N__45116),
            .I(N__45109));
    InMux I__10285 (
            .O(N__45115),
            .I(N__45109));
    InMux I__10284 (
            .O(N__45114),
            .I(N__45106));
    LocalMux I__10283 (
            .O(N__45109),
            .I(N__45103));
    LocalMux I__10282 (
            .O(N__45106),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv12 I__10281 (
            .O(N__45103),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__10280 (
            .O(N__45098),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__10279 (
            .O(N__45095),
            .I(N__45092));
    LocalMux I__10278 (
            .O(N__45092),
            .I(N__45089));
    Span4Mux_v I__10277 (
            .O(N__45089),
            .I(N__45086));
    Odrv4 I__10276 (
            .O(N__45086),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__10275 (
            .O(N__45083),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__10274 (
            .O(N__45080),
            .I(N__45077));
    LocalMux I__10273 (
            .O(N__45077),
            .I(N__45074));
    Odrv4 I__10272 (
            .O(N__45074),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__10271 (
            .O(N__45071),
            .I(bfn_17_20_0_));
    InMux I__10270 (
            .O(N__45068),
            .I(N__45065));
    LocalMux I__10269 (
            .O(N__45065),
            .I(N__45062));
    Odrv4 I__10268 (
            .O(N__45062),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__10267 (
            .O(N__45059),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__10266 (
            .O(N__45056),
            .I(N__45053));
    LocalMux I__10265 (
            .O(N__45053),
            .I(N__45050));
    Span4Mux_h I__10264 (
            .O(N__45050),
            .I(N__45047));
    Odrv4 I__10263 (
            .O(N__45047),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__10262 (
            .O(N__45044),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__10261 (
            .O(N__45041),
            .I(N__45038));
    LocalMux I__10260 (
            .O(N__45038),
            .I(N__45035));
    Odrv4 I__10259 (
            .O(N__45035),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__10258 (
            .O(N__45032),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__10257 (
            .O(N__45029),
            .I(N__45026));
    LocalMux I__10256 (
            .O(N__45026),
            .I(N__45023));
    Odrv4 I__10255 (
            .O(N__45023),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__10254 (
            .O(N__45020),
            .I(N__45015));
    InMux I__10253 (
            .O(N__45019),
            .I(N__45010));
    InMux I__10252 (
            .O(N__45018),
            .I(N__45010));
    LocalMux I__10251 (
            .O(N__45015),
            .I(N__45007));
    LocalMux I__10250 (
            .O(N__45010),
            .I(N__45004));
    Span4Mux_v I__10249 (
            .O(N__45007),
            .I(N__45001));
    Span4Mux_h I__10248 (
            .O(N__45004),
            .I(N__44998));
    Odrv4 I__10247 (
            .O(N__45001),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__10246 (
            .O(N__44998),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__10245 (
            .O(N__44993),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__10244 (
            .O(N__44990),
            .I(N__44987));
    LocalMux I__10243 (
            .O(N__44987),
            .I(N__44984));
    Span4Mux_h I__10242 (
            .O(N__44984),
            .I(N__44981));
    Odrv4 I__10241 (
            .O(N__44981),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__10240 (
            .O(N__44978),
            .I(N__44971));
    InMux I__10239 (
            .O(N__44977),
            .I(N__44971));
    InMux I__10238 (
            .O(N__44976),
            .I(N__44968));
    LocalMux I__10237 (
            .O(N__44971),
            .I(N__44965));
    LocalMux I__10236 (
            .O(N__44968),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__10235 (
            .O(N__44965),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__10234 (
            .O(N__44960),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    CascadeMux I__10233 (
            .O(N__44957),
            .I(N__44953));
    InMux I__10232 (
            .O(N__44956),
            .I(N__44950));
    InMux I__10231 (
            .O(N__44953),
            .I(N__44947));
    LocalMux I__10230 (
            .O(N__44950),
            .I(N__44944));
    LocalMux I__10229 (
            .O(N__44947),
            .I(N__44940));
    Span4Mux_h I__10228 (
            .O(N__44944),
            .I(N__44937));
    InMux I__10227 (
            .O(N__44943),
            .I(N__44934));
    Span4Mux_h I__10226 (
            .O(N__44940),
            .I(N__44931));
    Span4Mux_v I__10225 (
            .O(N__44937),
            .I(N__44928));
    LocalMux I__10224 (
            .O(N__44934),
            .I(N__44925));
    Odrv4 I__10223 (
            .O(N__44931),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__10222 (
            .O(N__44928),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv12 I__10221 (
            .O(N__44925),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__10220 (
            .O(N__44918),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__10219 (
            .O(N__44915),
            .I(N__44912));
    LocalMux I__10218 (
            .O(N__44912),
            .I(N__44909));
    Span4Mux_v I__10217 (
            .O(N__44909),
            .I(N__44906));
    Odrv4 I__10216 (
            .O(N__44906),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    CascadeMux I__10215 (
            .O(N__44903),
            .I(N__44899));
    InMux I__10214 (
            .O(N__44902),
            .I(N__44893));
    InMux I__10213 (
            .O(N__44899),
            .I(N__44893));
    InMux I__10212 (
            .O(N__44898),
            .I(N__44890));
    LocalMux I__10211 (
            .O(N__44893),
            .I(N__44887));
    LocalMux I__10210 (
            .O(N__44890),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__10209 (
            .O(N__44887),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__10208 (
            .O(N__44882),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__10207 (
            .O(N__44879),
            .I(N__44876));
    LocalMux I__10206 (
            .O(N__44876),
            .I(N__44873));
    Odrv4 I__10205 (
            .O(N__44873),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__10204 (
            .O(N__44870),
            .I(bfn_17_19_0_));
    InMux I__10203 (
            .O(N__44867),
            .I(N__44864));
    LocalMux I__10202 (
            .O(N__44864),
            .I(N__44861));
    Span4Mux_v I__10201 (
            .O(N__44861),
            .I(N__44858));
    Odrv4 I__10200 (
            .O(N__44858),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__10199 (
            .O(N__44855),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__10198 (
            .O(N__44852),
            .I(N__44849));
    LocalMux I__10197 (
            .O(N__44849),
            .I(N__44846));
    Span4Mux_h I__10196 (
            .O(N__44846),
            .I(N__44843));
    Span4Mux_v I__10195 (
            .O(N__44843),
            .I(N__44840));
    Odrv4 I__10194 (
            .O(N__44840),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__10193 (
            .O(N__44837),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__10192 (
            .O(N__44834),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__10191 (
            .O(N__44831),
            .I(N__44828));
    LocalMux I__10190 (
            .O(N__44828),
            .I(N__44825));
    Odrv4 I__10189 (
            .O(N__44825),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__10188 (
            .O(N__44822),
            .I(N__44818));
    InMux I__10187 (
            .O(N__44821),
            .I(N__44814));
    LocalMux I__10186 (
            .O(N__44818),
            .I(N__44811));
    InMux I__10185 (
            .O(N__44817),
            .I(N__44808));
    LocalMux I__10184 (
            .O(N__44814),
            .I(N__44805));
    Odrv4 I__10183 (
            .O(N__44811),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__10182 (
            .O(N__44808),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv12 I__10181 (
            .O(N__44805),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__10180 (
            .O(N__44798),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__10179 (
            .O(N__44795),
            .I(N__44789));
    InMux I__10178 (
            .O(N__44794),
            .I(N__44789));
    LocalMux I__10177 (
            .O(N__44789),
            .I(N__44785));
    InMux I__10176 (
            .O(N__44788),
            .I(N__44782));
    Span4Mux_v I__10175 (
            .O(N__44785),
            .I(N__44779));
    LocalMux I__10174 (
            .O(N__44782),
            .I(N__44776));
    Odrv4 I__10173 (
            .O(N__44779),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__10172 (
            .O(N__44776),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__10171 (
            .O(N__44771),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__10170 (
            .O(N__44768),
            .I(N__44765));
    LocalMux I__10169 (
            .O(N__44765),
            .I(N__44762));
    Odrv4 I__10168 (
            .O(N__44762),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__10167 (
            .O(N__44759),
            .I(N__44752));
    InMux I__10166 (
            .O(N__44758),
            .I(N__44752));
    InMux I__10165 (
            .O(N__44757),
            .I(N__44749));
    LocalMux I__10164 (
            .O(N__44752),
            .I(N__44746));
    LocalMux I__10163 (
            .O(N__44749),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv12 I__10162 (
            .O(N__44746),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__10161 (
            .O(N__44741),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__10160 (
            .O(N__44738),
            .I(N__44733));
    InMux I__10159 (
            .O(N__44737),
            .I(N__44730));
    InMux I__10158 (
            .O(N__44736),
            .I(N__44727));
    LocalMux I__10157 (
            .O(N__44733),
            .I(N__44724));
    LocalMux I__10156 (
            .O(N__44730),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__10155 (
            .O(N__44727),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__10154 (
            .O(N__44724),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__10153 (
            .O(N__44717),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__10152 (
            .O(N__44714),
            .I(N__44711));
    LocalMux I__10151 (
            .O(N__44711),
            .I(N__44708));
    Odrv4 I__10150 (
            .O(N__44708),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__10149 (
            .O(N__44705),
            .I(N__44698));
    InMux I__10148 (
            .O(N__44704),
            .I(N__44698));
    InMux I__10147 (
            .O(N__44703),
            .I(N__44695));
    LocalMux I__10146 (
            .O(N__44698),
            .I(N__44692));
    LocalMux I__10145 (
            .O(N__44695),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv4 I__10144 (
            .O(N__44692),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__10143 (
            .O(N__44687),
            .I(bfn_17_18_0_));
    InMux I__10142 (
            .O(N__44684),
            .I(N__44681));
    LocalMux I__10141 (
            .O(N__44681),
            .I(N__44678));
    Odrv4 I__10140 (
            .O(N__44678),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    CascadeMux I__10139 (
            .O(N__44675),
            .I(N__44672));
    InMux I__10138 (
            .O(N__44672),
            .I(N__44668));
    InMux I__10137 (
            .O(N__44671),
            .I(N__44665));
    LocalMux I__10136 (
            .O(N__44668),
            .I(N__44661));
    LocalMux I__10135 (
            .O(N__44665),
            .I(N__44658));
    InMux I__10134 (
            .O(N__44664),
            .I(N__44655));
    Span4Mux_h I__10133 (
            .O(N__44661),
            .I(N__44652));
    Span4Mux_h I__10132 (
            .O(N__44658),
            .I(N__44647));
    LocalMux I__10131 (
            .O(N__44655),
            .I(N__44647));
    Odrv4 I__10130 (
            .O(N__44652),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__10129 (
            .O(N__44647),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__10128 (
            .O(N__44642),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__10127 (
            .O(N__44639),
            .I(N__44636));
    LocalMux I__10126 (
            .O(N__44636),
            .I(N__44633));
    Span4Mux_h I__10125 (
            .O(N__44633),
            .I(N__44630));
    Odrv4 I__10124 (
            .O(N__44630),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__10123 (
            .O(N__44627),
            .I(N__44623));
    InMux I__10122 (
            .O(N__44626),
            .I(N__44619));
    LocalMux I__10121 (
            .O(N__44623),
            .I(N__44616));
    InMux I__10120 (
            .O(N__44622),
            .I(N__44613));
    LocalMux I__10119 (
            .O(N__44619),
            .I(N__44606));
    Span4Mux_h I__10118 (
            .O(N__44616),
            .I(N__44606));
    LocalMux I__10117 (
            .O(N__44613),
            .I(N__44606));
    Odrv4 I__10116 (
            .O(N__44606),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__10115 (
            .O(N__44603),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__10114 (
            .O(N__44600),
            .I(N__44597));
    LocalMux I__10113 (
            .O(N__44597),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__10112 (
            .O(N__44594),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    CascadeMux I__10111 (
            .O(N__44591),
            .I(N__44588));
    InMux I__10110 (
            .O(N__44588),
            .I(N__44585));
    LocalMux I__10109 (
            .O(N__44585),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    InMux I__10108 (
            .O(N__44582),
            .I(N__44579));
    LocalMux I__10107 (
            .O(N__44579),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    CascadeMux I__10106 (
            .O(N__44576),
            .I(N__44573));
    InMux I__10105 (
            .O(N__44573),
            .I(N__44568));
    InMux I__10104 (
            .O(N__44572),
            .I(N__44563));
    InMux I__10103 (
            .O(N__44571),
            .I(N__44563));
    LocalMux I__10102 (
            .O(N__44568),
            .I(N__44560));
    LocalMux I__10101 (
            .O(N__44563),
            .I(N__44557));
    Span4Mux_h I__10100 (
            .O(N__44560),
            .I(N__44553));
    Span12Mux_s10_h I__10099 (
            .O(N__44557),
            .I(N__44550));
    InMux I__10098 (
            .O(N__44556),
            .I(N__44547));
    Odrv4 I__10097 (
            .O(N__44553),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv12 I__10096 (
            .O(N__44550),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__10095 (
            .O(N__44547),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    CascadeMux I__10094 (
            .O(N__44540),
            .I(N__44537));
    InMux I__10093 (
            .O(N__44537),
            .I(N__44532));
    InMux I__10092 (
            .O(N__44536),
            .I(N__44529));
    InMux I__10091 (
            .O(N__44535),
            .I(N__44526));
    LocalMux I__10090 (
            .O(N__44532),
            .I(N__44523));
    LocalMux I__10089 (
            .O(N__44529),
            .I(N__44520));
    LocalMux I__10088 (
            .O(N__44526),
            .I(N__44517));
    Span4Mux_h I__10087 (
            .O(N__44523),
            .I(N__44514));
    Span4Mux_h I__10086 (
            .O(N__44520),
            .I(N__44511));
    Span4Mux_h I__10085 (
            .O(N__44517),
            .I(N__44508));
    Span4Mux_v I__10084 (
            .O(N__44514),
            .I(N__44504));
    Span4Mux_v I__10083 (
            .O(N__44511),
            .I(N__44501));
    Span4Mux_v I__10082 (
            .O(N__44508),
            .I(N__44498));
    InMux I__10081 (
            .O(N__44507),
            .I(N__44495));
    Odrv4 I__10080 (
            .O(N__44504),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10079 (
            .O(N__44501),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10078 (
            .O(N__44498),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__10077 (
            .O(N__44495),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10076 (
            .O(N__44486),
            .I(N__44483));
    LocalMux I__10075 (
            .O(N__44483),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    InMux I__10074 (
            .O(N__44480),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__10073 (
            .O(N__44477),
            .I(N__44474));
    LocalMux I__10072 (
            .O(N__44474),
            .I(N__44471));
    Span4Mux_h I__10071 (
            .O(N__44471),
            .I(N__44468));
    Odrv4 I__10070 (
            .O(N__44468),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__10069 (
            .O(N__44465),
            .I(N__44462));
    LocalMux I__10068 (
            .O(N__44462),
            .I(N__44457));
    InMux I__10067 (
            .O(N__44461),
            .I(N__44452));
    InMux I__10066 (
            .O(N__44460),
            .I(N__44452));
    Span4Mux_v I__10065 (
            .O(N__44457),
            .I(N__44449));
    LocalMux I__10064 (
            .O(N__44452),
            .I(N__44446));
    Odrv4 I__10063 (
            .O(N__44449),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__10062 (
            .O(N__44446),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__10061 (
            .O(N__44441),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__10060 (
            .O(N__44438),
            .I(N__44435));
    LocalMux I__10059 (
            .O(N__44435),
            .I(N__44432));
    Span4Mux_h I__10058 (
            .O(N__44432),
            .I(N__44429));
    Odrv4 I__10057 (
            .O(N__44429),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__10056 (
            .O(N__44426),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__10055 (
            .O(N__44423),
            .I(N__44420));
    LocalMux I__10054 (
            .O(N__44420),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    InMux I__10053 (
            .O(N__44417),
            .I(N__44413));
    InMux I__10052 (
            .O(N__44416),
            .I(N__44409));
    LocalMux I__10051 (
            .O(N__44413),
            .I(N__44406));
    InMux I__10050 (
            .O(N__44412),
            .I(N__44403));
    LocalMux I__10049 (
            .O(N__44409),
            .I(N__44400));
    Span4Mux_h I__10048 (
            .O(N__44406),
            .I(N__44397));
    LocalMux I__10047 (
            .O(N__44403),
            .I(N__44393));
    Span4Mux_h I__10046 (
            .O(N__44400),
            .I(N__44388));
    Span4Mux_v I__10045 (
            .O(N__44397),
            .I(N__44388));
    InMux I__10044 (
            .O(N__44396),
            .I(N__44385));
    Odrv12 I__10043 (
            .O(N__44393),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__10042 (
            .O(N__44388),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__10041 (
            .O(N__44385),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    CascadeMux I__10040 (
            .O(N__44378),
            .I(N__44373));
    InMux I__10039 (
            .O(N__44377),
            .I(N__44368));
    InMux I__10038 (
            .O(N__44376),
            .I(N__44368));
    InMux I__10037 (
            .O(N__44373),
            .I(N__44365));
    LocalMux I__10036 (
            .O(N__44368),
            .I(N__44362));
    LocalMux I__10035 (
            .O(N__44365),
            .I(N__44359));
    Span4Mux_h I__10034 (
            .O(N__44362),
            .I(N__44356));
    Span4Mux_h I__10033 (
            .O(N__44359),
            .I(N__44352));
    Span4Mux_v I__10032 (
            .O(N__44356),
            .I(N__44349));
    InMux I__10031 (
            .O(N__44355),
            .I(N__44346));
    Odrv4 I__10030 (
            .O(N__44352),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__10029 (
            .O(N__44349),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__10028 (
            .O(N__44346),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    CascadeMux I__10027 (
            .O(N__44339),
            .I(N__44336));
    InMux I__10026 (
            .O(N__44336),
            .I(N__44329));
    InMux I__10025 (
            .O(N__44335),
            .I(N__44329));
    InMux I__10024 (
            .O(N__44334),
            .I(N__44326));
    LocalMux I__10023 (
            .O(N__44329),
            .I(N__44323));
    LocalMux I__10022 (
            .O(N__44326),
            .I(N__44318));
    Span4Mux_v I__10021 (
            .O(N__44323),
            .I(N__44318));
    Span4Mux_v I__10020 (
            .O(N__44318),
            .I(N__44314));
    InMux I__10019 (
            .O(N__44317),
            .I(N__44311));
    Odrv4 I__10018 (
            .O(N__44314),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__10017 (
            .O(N__44311),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    CascadeMux I__10016 (
            .O(N__44306),
            .I(N__44303));
    InMux I__10015 (
            .O(N__44303),
            .I(N__44300));
    LocalMux I__10014 (
            .O(N__44300),
            .I(N__44297));
    Odrv4 I__10013 (
            .O(N__44297),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    InMux I__10012 (
            .O(N__44294),
            .I(N__44291));
    LocalMux I__10011 (
            .O(N__44291),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    CascadeMux I__10010 (
            .O(N__44288),
            .I(N__44285));
    InMux I__10009 (
            .O(N__44285),
            .I(N__44282));
    LocalMux I__10008 (
            .O(N__44282),
            .I(N__44279));
    Odrv4 I__10007 (
            .O(N__44279),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    CascadeMux I__10006 (
            .O(N__44276),
            .I(N__44273));
    InMux I__10005 (
            .O(N__44273),
            .I(N__44270));
    LocalMux I__10004 (
            .O(N__44270),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    CascadeMux I__10003 (
            .O(N__44267),
            .I(N__44264));
    InMux I__10002 (
            .O(N__44264),
            .I(N__44259));
    InMux I__10001 (
            .O(N__44263),
            .I(N__44256));
    InMux I__10000 (
            .O(N__44262),
            .I(N__44253));
    LocalMux I__9999 (
            .O(N__44259),
            .I(N__44250));
    LocalMux I__9998 (
            .O(N__44256),
            .I(N__44247));
    LocalMux I__9997 (
            .O(N__44253),
            .I(N__44244));
    Span4Mux_h I__9996 (
            .O(N__44250),
            .I(N__44241));
    Span4Mux_h I__9995 (
            .O(N__44247),
            .I(N__44238));
    Span4Mux_h I__9994 (
            .O(N__44244),
            .I(N__44232));
    Span4Mux_v I__9993 (
            .O(N__44241),
            .I(N__44232));
    Span4Mux_v I__9992 (
            .O(N__44238),
            .I(N__44229));
    InMux I__9991 (
            .O(N__44237),
            .I(N__44226));
    Odrv4 I__9990 (
            .O(N__44232),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__9989 (
            .O(N__44229),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__9988 (
            .O(N__44226),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    CascadeMux I__9987 (
            .O(N__44219),
            .I(N__44216));
    InMux I__9986 (
            .O(N__44216),
            .I(N__44213));
    LocalMux I__9985 (
            .O(N__44213),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    CascadeMux I__9984 (
            .O(N__44210),
            .I(N__44207));
    InMux I__9983 (
            .O(N__44207),
            .I(N__44200));
    InMux I__9982 (
            .O(N__44206),
            .I(N__44200));
    InMux I__9981 (
            .O(N__44205),
            .I(N__44197));
    LocalMux I__9980 (
            .O(N__44200),
            .I(N__44194));
    LocalMux I__9979 (
            .O(N__44197),
            .I(N__44190));
    Span12Mux_s10_h I__9978 (
            .O(N__44194),
            .I(N__44187));
    InMux I__9977 (
            .O(N__44193),
            .I(N__44184));
    Odrv4 I__9976 (
            .O(N__44190),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv12 I__9975 (
            .O(N__44187),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__9974 (
            .O(N__44184),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__9973 (
            .O(N__44177),
            .I(N__44174));
    LocalMux I__9972 (
            .O(N__44174),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__9971 (
            .O(N__44171),
            .I(N__44168));
    InMux I__9970 (
            .O(N__44168),
            .I(N__44162));
    InMux I__9969 (
            .O(N__44167),
            .I(N__44162));
    LocalMux I__9968 (
            .O(N__44162),
            .I(N__44158));
    InMux I__9967 (
            .O(N__44161),
            .I(N__44155));
    Span4Mux_h I__9966 (
            .O(N__44158),
            .I(N__44152));
    LocalMux I__9965 (
            .O(N__44155),
            .I(N__44146));
    Span4Mux_v I__9964 (
            .O(N__44152),
            .I(N__44146));
    InMux I__9963 (
            .O(N__44151),
            .I(N__44143));
    Odrv4 I__9962 (
            .O(N__44146),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__9961 (
            .O(N__44143),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    CascadeMux I__9960 (
            .O(N__44138),
            .I(N__44135));
    InMux I__9959 (
            .O(N__44135),
            .I(N__44132));
    LocalMux I__9958 (
            .O(N__44132),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    CascadeMux I__9957 (
            .O(N__44129),
            .I(N__44126));
    InMux I__9956 (
            .O(N__44126),
            .I(N__44123));
    LocalMux I__9955 (
            .O(N__44123),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    InMux I__9954 (
            .O(N__44120),
            .I(N__44104));
    InMux I__9953 (
            .O(N__44119),
            .I(N__44104));
    InMux I__9952 (
            .O(N__44118),
            .I(N__44104));
    InMux I__9951 (
            .O(N__44117),
            .I(N__44104));
    InMux I__9950 (
            .O(N__44116),
            .I(N__44095));
    InMux I__9949 (
            .O(N__44115),
            .I(N__44095));
    InMux I__9948 (
            .O(N__44114),
            .I(N__44095));
    InMux I__9947 (
            .O(N__44113),
            .I(N__44095));
    LocalMux I__9946 (
            .O(N__44104),
            .I(N__44072));
    LocalMux I__9945 (
            .O(N__44095),
            .I(N__44072));
    InMux I__9944 (
            .O(N__44094),
            .I(N__44063));
    InMux I__9943 (
            .O(N__44093),
            .I(N__44063));
    InMux I__9942 (
            .O(N__44092),
            .I(N__44063));
    InMux I__9941 (
            .O(N__44091),
            .I(N__44063));
    InMux I__9940 (
            .O(N__44090),
            .I(N__44058));
    InMux I__9939 (
            .O(N__44089),
            .I(N__44058));
    InMux I__9938 (
            .O(N__44088),
            .I(N__44045));
    InMux I__9937 (
            .O(N__44087),
            .I(N__44045));
    InMux I__9936 (
            .O(N__44086),
            .I(N__44045));
    InMux I__9935 (
            .O(N__44085),
            .I(N__44045));
    InMux I__9934 (
            .O(N__44084),
            .I(N__44036));
    InMux I__9933 (
            .O(N__44083),
            .I(N__44036));
    InMux I__9932 (
            .O(N__44082),
            .I(N__44036));
    InMux I__9931 (
            .O(N__44081),
            .I(N__44036));
    InMux I__9930 (
            .O(N__44080),
            .I(N__44027));
    InMux I__9929 (
            .O(N__44079),
            .I(N__44027));
    InMux I__9928 (
            .O(N__44078),
            .I(N__44027));
    InMux I__9927 (
            .O(N__44077),
            .I(N__44027));
    Span4Mux_v I__9926 (
            .O(N__44072),
            .I(N__44020));
    LocalMux I__9925 (
            .O(N__44063),
            .I(N__44020));
    LocalMux I__9924 (
            .O(N__44058),
            .I(N__44020));
    InMux I__9923 (
            .O(N__44057),
            .I(N__44011));
    InMux I__9922 (
            .O(N__44056),
            .I(N__44011));
    InMux I__9921 (
            .O(N__44055),
            .I(N__44011));
    InMux I__9920 (
            .O(N__44054),
            .I(N__44011));
    LocalMux I__9919 (
            .O(N__44045),
            .I(N__44006));
    LocalMux I__9918 (
            .O(N__44036),
            .I(N__44006));
    LocalMux I__9917 (
            .O(N__44027),
            .I(N__44001));
    Span4Mux_v I__9916 (
            .O(N__44020),
            .I(N__44001));
    LocalMux I__9915 (
            .O(N__44011),
            .I(N__43998));
    Span4Mux_v I__9914 (
            .O(N__44006),
            .I(N__43993));
    Span4Mux_h I__9913 (
            .O(N__44001),
            .I(N__43993));
    Odrv4 I__9912 (
            .O(N__43998),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9911 (
            .O(N__43993),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9910 (
            .O(N__43988),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__9909 (
            .O(N__43985),
            .I(N__43981));
    InMux I__9908 (
            .O(N__43984),
            .I(N__43978));
    LocalMux I__9907 (
            .O(N__43981),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__9906 (
            .O(N__43978),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__9905 (
            .O(N__43973),
            .I(N__43970));
    LocalMux I__9904 (
            .O(N__43970),
            .I(N__43966));
    CEMux I__9903 (
            .O(N__43969),
            .I(N__43962));
    Span4Mux_v I__9902 (
            .O(N__43966),
            .I(N__43959));
    CEMux I__9901 (
            .O(N__43965),
            .I(N__43956));
    LocalMux I__9900 (
            .O(N__43962),
            .I(N__43948));
    Span4Mux_h I__9899 (
            .O(N__43959),
            .I(N__43948));
    LocalMux I__9898 (
            .O(N__43956),
            .I(N__43948));
    CEMux I__9897 (
            .O(N__43955),
            .I(N__43945));
    Sp12to4 I__9896 (
            .O(N__43948),
            .I(N__43940));
    LocalMux I__9895 (
            .O(N__43945),
            .I(N__43940));
    Odrv12 I__9894 (
            .O(N__43940),
            .I(\delay_measurement_inst.delay_tr_timer.N_305_i ));
    InMux I__9893 (
            .O(N__43937),
            .I(N__43934));
    LocalMux I__9892 (
            .O(N__43934),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__9891 (
            .O(N__43931),
            .I(N__43927));
    InMux I__9890 (
            .O(N__43930),
            .I(N__43924));
    LocalMux I__9889 (
            .O(N__43927),
            .I(N__43921));
    LocalMux I__9888 (
            .O(N__43924),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv12 I__9887 (
            .O(N__43921),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__9886 (
            .O(N__43916),
            .I(N__43911));
    InMux I__9885 (
            .O(N__43915),
            .I(N__43908));
    InMux I__9884 (
            .O(N__43914),
            .I(N__43905));
    LocalMux I__9883 (
            .O(N__43911),
            .I(N__43900));
    LocalMux I__9882 (
            .O(N__43908),
            .I(N__43900));
    LocalMux I__9881 (
            .O(N__43905),
            .I(N__43895));
    Span4Mux_v I__9880 (
            .O(N__43900),
            .I(N__43895));
    Odrv4 I__9879 (
            .O(N__43895),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    CascadeMux I__9878 (
            .O(N__43892),
            .I(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ));
    InMux I__9877 (
            .O(N__43889),
            .I(N__43886));
    LocalMux I__9876 (
            .O(N__43886),
            .I(N__43883));
    Span4Mux_h I__9875 (
            .O(N__43883),
            .I(N__43875));
    InMux I__9874 (
            .O(N__43882),
            .I(N__43872));
    InMux I__9873 (
            .O(N__43881),
            .I(N__43863));
    InMux I__9872 (
            .O(N__43880),
            .I(N__43863));
    InMux I__9871 (
            .O(N__43879),
            .I(N__43863));
    InMux I__9870 (
            .O(N__43878),
            .I(N__43863));
    Odrv4 I__9869 (
            .O(N__43875),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9868 (
            .O(N__43872),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9867 (
            .O(N__43863),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__9866 (
            .O(N__43856),
            .I(N__43852));
    InMux I__9865 (
            .O(N__43855),
            .I(N__43849));
    LocalMux I__9864 (
            .O(N__43852),
            .I(N__43846));
    LocalMux I__9863 (
            .O(N__43849),
            .I(N__43843));
    Span4Mux_h I__9862 (
            .O(N__43846),
            .I(N__43840));
    Span4Mux_h I__9861 (
            .O(N__43843),
            .I(N__43837));
    Span4Mux_v I__9860 (
            .O(N__43840),
            .I(N__43834));
    Span4Mux_h I__9859 (
            .O(N__43837),
            .I(N__43831));
    Odrv4 I__9858 (
            .O(N__43834),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    Odrv4 I__9857 (
            .O(N__43831),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    InMux I__9856 (
            .O(N__43826),
            .I(N__43808));
    InMux I__9855 (
            .O(N__43825),
            .I(N__43808));
    InMux I__9854 (
            .O(N__43824),
            .I(N__43808));
    CascadeMux I__9853 (
            .O(N__43823),
            .I(N__43805));
    CascadeMux I__9852 (
            .O(N__43822),
            .I(N__43801));
    InMux I__9851 (
            .O(N__43821),
            .I(N__43779));
    InMux I__9850 (
            .O(N__43820),
            .I(N__43779));
    InMux I__9849 (
            .O(N__43819),
            .I(N__43779));
    InMux I__9848 (
            .O(N__43818),
            .I(N__43779));
    InMux I__9847 (
            .O(N__43817),
            .I(N__43779));
    InMux I__9846 (
            .O(N__43816),
            .I(N__43779));
    InMux I__9845 (
            .O(N__43815),
            .I(N__43779));
    LocalMux I__9844 (
            .O(N__43808),
            .I(N__43772));
    InMux I__9843 (
            .O(N__43805),
            .I(N__43767));
    InMux I__9842 (
            .O(N__43804),
            .I(N__43767));
    InMux I__9841 (
            .O(N__43801),
            .I(N__43750));
    InMux I__9840 (
            .O(N__43800),
            .I(N__43750));
    InMux I__9839 (
            .O(N__43799),
            .I(N__43750));
    InMux I__9838 (
            .O(N__43798),
            .I(N__43750));
    InMux I__9837 (
            .O(N__43797),
            .I(N__43750));
    InMux I__9836 (
            .O(N__43796),
            .I(N__43750));
    InMux I__9835 (
            .O(N__43795),
            .I(N__43750));
    InMux I__9834 (
            .O(N__43794),
            .I(N__43750));
    LocalMux I__9833 (
            .O(N__43779),
            .I(N__43747));
    InMux I__9832 (
            .O(N__43778),
            .I(N__43738));
    InMux I__9831 (
            .O(N__43777),
            .I(N__43738));
    InMux I__9830 (
            .O(N__43776),
            .I(N__43738));
    InMux I__9829 (
            .O(N__43775),
            .I(N__43738));
    Span4Mux_v I__9828 (
            .O(N__43772),
            .I(N__43735));
    LocalMux I__9827 (
            .O(N__43767),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__9826 (
            .O(N__43750),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__9825 (
            .O(N__43747),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__9824 (
            .O(N__43738),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__9823 (
            .O(N__43735),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__9822 (
            .O(N__43724),
            .I(N__43713));
    CascadeMux I__9821 (
            .O(N__43723),
            .I(N__43709));
    CascadeMux I__9820 (
            .O(N__43722),
            .I(N__43705));
    CascadeMux I__9819 (
            .O(N__43721),
            .I(N__43701));
    CascadeMux I__9818 (
            .O(N__43720),
            .I(N__43697));
    CascadeMux I__9817 (
            .O(N__43719),
            .I(N__43692));
    CascadeMux I__9816 (
            .O(N__43718),
            .I(N__43688));
    CascadeMux I__9815 (
            .O(N__43717),
            .I(N__43684));
    InMux I__9814 (
            .O(N__43716),
            .I(N__43678));
    InMux I__9813 (
            .O(N__43713),
            .I(N__43678));
    InMux I__9812 (
            .O(N__43712),
            .I(N__43661));
    InMux I__9811 (
            .O(N__43709),
            .I(N__43661));
    InMux I__9810 (
            .O(N__43708),
            .I(N__43661));
    InMux I__9809 (
            .O(N__43705),
            .I(N__43661));
    InMux I__9808 (
            .O(N__43704),
            .I(N__43661));
    InMux I__9807 (
            .O(N__43701),
            .I(N__43661));
    InMux I__9806 (
            .O(N__43700),
            .I(N__43661));
    InMux I__9805 (
            .O(N__43697),
            .I(N__43661));
    InMux I__9804 (
            .O(N__43696),
            .I(N__43657));
    InMux I__9803 (
            .O(N__43695),
            .I(N__43644));
    InMux I__9802 (
            .O(N__43692),
            .I(N__43644));
    InMux I__9801 (
            .O(N__43691),
            .I(N__43644));
    InMux I__9800 (
            .O(N__43688),
            .I(N__43644));
    InMux I__9799 (
            .O(N__43687),
            .I(N__43644));
    InMux I__9798 (
            .O(N__43684),
            .I(N__43644));
    CascadeMux I__9797 (
            .O(N__43683),
            .I(N__43641));
    LocalMux I__9796 (
            .O(N__43678),
            .I(N__43635));
    LocalMux I__9795 (
            .O(N__43661),
            .I(N__43635));
    CascadeMux I__9794 (
            .O(N__43660),
            .I(N__43631));
    LocalMux I__9793 (
            .O(N__43657),
            .I(N__43624));
    LocalMux I__9792 (
            .O(N__43644),
            .I(N__43624));
    InMux I__9791 (
            .O(N__43641),
            .I(N__43619));
    InMux I__9790 (
            .O(N__43640),
            .I(N__43619));
    Span4Mux_v I__9789 (
            .O(N__43635),
            .I(N__43616));
    InMux I__9788 (
            .O(N__43634),
            .I(N__43607));
    InMux I__9787 (
            .O(N__43631),
            .I(N__43607));
    InMux I__9786 (
            .O(N__43630),
            .I(N__43607));
    InMux I__9785 (
            .O(N__43629),
            .I(N__43607));
    Span4Mux_h I__9784 (
            .O(N__43624),
            .I(N__43602));
    LocalMux I__9783 (
            .O(N__43619),
            .I(N__43602));
    Sp12to4 I__9782 (
            .O(N__43616),
            .I(N__43596));
    LocalMux I__9781 (
            .O(N__43607),
            .I(N__43596));
    Span4Mux_v I__9780 (
            .O(N__43602),
            .I(N__43593));
    InMux I__9779 (
            .O(N__43601),
            .I(N__43590));
    Span12Mux_h I__9778 (
            .O(N__43596),
            .I(N__43587));
    Span4Mux_h I__9777 (
            .O(N__43593),
            .I(N__43584));
    LocalMux I__9776 (
            .O(N__43590),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__9775 (
            .O(N__43587),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__9774 (
            .O(N__43584),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__9773 (
            .O(N__43577),
            .I(N__43572));
    CascadeMux I__9772 (
            .O(N__43576),
            .I(N__43569));
    CascadeMux I__9771 (
            .O(N__43575),
            .I(N__43566));
    InMux I__9770 (
            .O(N__43572),
            .I(N__43547));
    InMux I__9769 (
            .O(N__43569),
            .I(N__43547));
    InMux I__9768 (
            .O(N__43566),
            .I(N__43547));
    InMux I__9767 (
            .O(N__43565),
            .I(N__43538));
    InMux I__9766 (
            .O(N__43564),
            .I(N__43538));
    InMux I__9765 (
            .O(N__43563),
            .I(N__43538));
    InMux I__9764 (
            .O(N__43562),
            .I(N__43538));
    InMux I__9763 (
            .O(N__43561),
            .I(N__43533));
    InMux I__9762 (
            .O(N__43560),
            .I(N__43533));
    InMux I__9761 (
            .O(N__43559),
            .I(N__43530));
    CascadeMux I__9760 (
            .O(N__43558),
            .I(N__43527));
    CascadeMux I__9759 (
            .O(N__43557),
            .I(N__43523));
    CascadeMux I__9758 (
            .O(N__43556),
            .I(N__43520));
    CascadeMux I__9757 (
            .O(N__43555),
            .I(N__43510));
    CascadeMux I__9756 (
            .O(N__43554),
            .I(N__43507));
    LocalMux I__9755 (
            .O(N__43547),
            .I(N__43497));
    LocalMux I__9754 (
            .O(N__43538),
            .I(N__43497));
    LocalMux I__9753 (
            .O(N__43533),
            .I(N__43497));
    LocalMux I__9752 (
            .O(N__43530),
            .I(N__43497));
    InMux I__9751 (
            .O(N__43527),
            .I(N__43488));
    InMux I__9750 (
            .O(N__43526),
            .I(N__43488));
    InMux I__9749 (
            .O(N__43523),
            .I(N__43488));
    InMux I__9748 (
            .O(N__43520),
            .I(N__43488));
    InMux I__9747 (
            .O(N__43519),
            .I(N__43483));
    InMux I__9746 (
            .O(N__43518),
            .I(N__43483));
    InMux I__9745 (
            .O(N__43517),
            .I(N__43480));
    InMux I__9744 (
            .O(N__43516),
            .I(N__43471));
    InMux I__9743 (
            .O(N__43515),
            .I(N__43471));
    InMux I__9742 (
            .O(N__43514),
            .I(N__43471));
    InMux I__9741 (
            .O(N__43513),
            .I(N__43471));
    InMux I__9740 (
            .O(N__43510),
            .I(N__43464));
    InMux I__9739 (
            .O(N__43507),
            .I(N__43464));
    InMux I__9738 (
            .O(N__43506),
            .I(N__43464));
    Span4Mux_h I__9737 (
            .O(N__43497),
            .I(N__43461));
    LocalMux I__9736 (
            .O(N__43488),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__9735 (
            .O(N__43483),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__9734 (
            .O(N__43480),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__9733 (
            .O(N__43471),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__9732 (
            .O(N__43464),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__9731 (
            .O(N__43461),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__9730 (
            .O(N__43448),
            .I(N__43445));
    LocalMux I__9729 (
            .O(N__43445),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__9728 (
            .O(N__43442),
            .I(N__43439));
    LocalMux I__9727 (
            .O(N__43439),
            .I(N__43436));
    Span4Mux_v I__9726 (
            .O(N__43436),
            .I(N__43432));
    InMux I__9725 (
            .O(N__43435),
            .I(N__43429));
    Span4Mux_v I__9724 (
            .O(N__43432),
            .I(N__43426));
    LocalMux I__9723 (
            .O(N__43429),
            .I(N__43423));
    Span4Mux_v I__9722 (
            .O(N__43426),
            .I(N__43420));
    Span12Mux_h I__9721 (
            .O(N__43423),
            .I(N__43416));
    Span4Mux_v I__9720 (
            .O(N__43420),
            .I(N__43413));
    InMux I__9719 (
            .O(N__43419),
            .I(N__43410));
    Odrv12 I__9718 (
            .O(N__43416),
            .I(il_min_comp1_D2));
    Odrv4 I__9717 (
            .O(N__43413),
            .I(il_min_comp1_D2));
    LocalMux I__9716 (
            .O(N__43410),
            .I(il_min_comp1_D2));
    InMux I__9715 (
            .O(N__43403),
            .I(N__43398));
    InMux I__9714 (
            .O(N__43402),
            .I(N__43393));
    InMux I__9713 (
            .O(N__43401),
            .I(N__43393));
    LocalMux I__9712 (
            .O(N__43398),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__9711 (
            .O(N__43393),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__9710 (
            .O(N__43388),
            .I(N__43385));
    InMux I__9709 (
            .O(N__43385),
            .I(N__43382));
    LocalMux I__9708 (
            .O(N__43382),
            .I(N__43377));
    InMux I__9707 (
            .O(N__43381),
            .I(N__43374));
    InMux I__9706 (
            .O(N__43380),
            .I(N__43371));
    Span4Mux_v I__9705 (
            .O(N__43377),
            .I(N__43368));
    LocalMux I__9704 (
            .O(N__43374),
            .I(N__43364));
    LocalMux I__9703 (
            .O(N__43371),
            .I(N__43361));
    Span4Mux_v I__9702 (
            .O(N__43368),
            .I(N__43358));
    CascadeMux I__9701 (
            .O(N__43367),
            .I(N__43355));
    Span12Mux_s7_v I__9700 (
            .O(N__43364),
            .I(N__43352));
    Span4Mux_v I__9699 (
            .O(N__43361),
            .I(N__43347));
    Span4Mux_h I__9698 (
            .O(N__43358),
            .I(N__43347));
    InMux I__9697 (
            .O(N__43355),
            .I(N__43344));
    Span12Mux_v I__9696 (
            .O(N__43352),
            .I(N__43341));
    Odrv4 I__9695 (
            .O(N__43347),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__9694 (
            .O(N__43344),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__9693 (
            .O(N__43341),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__9692 (
            .O(N__43334),
            .I(N__43330));
    InMux I__9691 (
            .O(N__43333),
            .I(N__43327));
    LocalMux I__9690 (
            .O(N__43330),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__9689 (
            .O(N__43327),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__9688 (
            .O(N__43322),
            .I(N__43317));
    InMux I__9687 (
            .O(N__43321),
            .I(N__43312));
    InMux I__9686 (
            .O(N__43320),
            .I(N__43312));
    LocalMux I__9685 (
            .O(N__43317),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__9684 (
            .O(N__43312),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__9683 (
            .O(N__43307),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__9682 (
            .O(N__43304),
            .I(N__43299));
    InMux I__9681 (
            .O(N__43303),
            .I(N__43294));
    InMux I__9680 (
            .O(N__43302),
            .I(N__43294));
    LocalMux I__9679 (
            .O(N__43299),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__9678 (
            .O(N__43294),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__9677 (
            .O(N__43289),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__9676 (
            .O(N__43286),
            .I(N__43281));
    CascadeMux I__9675 (
            .O(N__43285),
            .I(N__43278));
    InMux I__9674 (
            .O(N__43284),
            .I(N__43275));
    InMux I__9673 (
            .O(N__43281),
            .I(N__43270));
    InMux I__9672 (
            .O(N__43278),
            .I(N__43270));
    LocalMux I__9671 (
            .O(N__43275),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__9670 (
            .O(N__43270),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__9669 (
            .O(N__43265),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__9668 (
            .O(N__43262),
            .I(N__43257));
    CascadeMux I__9667 (
            .O(N__43261),
            .I(N__43254));
    InMux I__9666 (
            .O(N__43260),
            .I(N__43251));
    InMux I__9665 (
            .O(N__43257),
            .I(N__43246));
    InMux I__9664 (
            .O(N__43254),
            .I(N__43246));
    LocalMux I__9663 (
            .O(N__43251),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__9662 (
            .O(N__43246),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__9661 (
            .O(N__43241),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9660 (
            .O(N__43238),
            .I(N__43233));
    InMux I__9659 (
            .O(N__43237),
            .I(N__43230));
    InMux I__9658 (
            .O(N__43236),
            .I(N__43227));
    LocalMux I__9657 (
            .O(N__43233),
            .I(N__43224));
    LocalMux I__9656 (
            .O(N__43230),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__9655 (
            .O(N__43227),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__9654 (
            .O(N__43224),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__9653 (
            .O(N__43217),
            .I(bfn_17_10_0_));
    InMux I__9652 (
            .O(N__43214),
            .I(N__43209));
    InMux I__9651 (
            .O(N__43213),
            .I(N__43206));
    InMux I__9650 (
            .O(N__43212),
            .I(N__43203));
    LocalMux I__9649 (
            .O(N__43209),
            .I(N__43200));
    LocalMux I__9648 (
            .O(N__43206),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__9647 (
            .O(N__43203),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__9646 (
            .O(N__43200),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__9645 (
            .O(N__43193),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__9644 (
            .O(N__43190),
            .I(N__43185));
    CascadeMux I__9643 (
            .O(N__43189),
            .I(N__43182));
    InMux I__9642 (
            .O(N__43188),
            .I(N__43179));
    InMux I__9641 (
            .O(N__43185),
            .I(N__43174));
    InMux I__9640 (
            .O(N__43182),
            .I(N__43174));
    LocalMux I__9639 (
            .O(N__43179),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__9638 (
            .O(N__43174),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__9637 (
            .O(N__43169),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__9636 (
            .O(N__43166),
            .I(N__43161));
    CascadeMux I__9635 (
            .O(N__43165),
            .I(N__43158));
    InMux I__9634 (
            .O(N__43164),
            .I(N__43155));
    InMux I__9633 (
            .O(N__43161),
            .I(N__43150));
    InMux I__9632 (
            .O(N__43158),
            .I(N__43150));
    LocalMux I__9631 (
            .O(N__43155),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__9630 (
            .O(N__43150),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__9629 (
            .O(N__43145),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9628 (
            .O(N__43142),
            .I(N__43138));
    InMux I__9627 (
            .O(N__43141),
            .I(N__43135));
    LocalMux I__9626 (
            .O(N__43138),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__9625 (
            .O(N__43135),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__9624 (
            .O(N__43130),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__9623 (
            .O(N__43127),
            .I(N__43122));
    InMux I__9622 (
            .O(N__43126),
            .I(N__43117));
    InMux I__9621 (
            .O(N__43125),
            .I(N__43117));
    LocalMux I__9620 (
            .O(N__43122),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__9619 (
            .O(N__43117),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__9618 (
            .O(N__43112),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__9617 (
            .O(N__43109),
            .I(N__43104));
    InMux I__9616 (
            .O(N__43108),
            .I(N__43099));
    InMux I__9615 (
            .O(N__43107),
            .I(N__43099));
    LocalMux I__9614 (
            .O(N__43104),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__9613 (
            .O(N__43099),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__9612 (
            .O(N__43094),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__9611 (
            .O(N__43091),
            .I(N__43086));
    CascadeMux I__9610 (
            .O(N__43090),
            .I(N__43083));
    InMux I__9609 (
            .O(N__43089),
            .I(N__43080));
    InMux I__9608 (
            .O(N__43086),
            .I(N__43075));
    InMux I__9607 (
            .O(N__43083),
            .I(N__43075));
    LocalMux I__9606 (
            .O(N__43080),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__9605 (
            .O(N__43075),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__9604 (
            .O(N__43070),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__9603 (
            .O(N__43067),
            .I(N__43062));
    CascadeMux I__9602 (
            .O(N__43066),
            .I(N__43059));
    InMux I__9601 (
            .O(N__43065),
            .I(N__43056));
    InMux I__9600 (
            .O(N__43062),
            .I(N__43051));
    InMux I__9599 (
            .O(N__43059),
            .I(N__43051));
    LocalMux I__9598 (
            .O(N__43056),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__9597 (
            .O(N__43051),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__9596 (
            .O(N__43046),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__9595 (
            .O(N__43043),
            .I(N__43038));
    InMux I__9594 (
            .O(N__43042),
            .I(N__43035));
    InMux I__9593 (
            .O(N__43041),
            .I(N__43032));
    LocalMux I__9592 (
            .O(N__43038),
            .I(N__43029));
    LocalMux I__9591 (
            .O(N__43035),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__9590 (
            .O(N__43032),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__9589 (
            .O(N__43029),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__9588 (
            .O(N__43022),
            .I(bfn_17_9_0_));
    InMux I__9587 (
            .O(N__43019),
            .I(N__43014));
    InMux I__9586 (
            .O(N__43018),
            .I(N__43011));
    InMux I__9585 (
            .O(N__43017),
            .I(N__43008));
    LocalMux I__9584 (
            .O(N__43014),
            .I(N__43005));
    LocalMux I__9583 (
            .O(N__43011),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__9582 (
            .O(N__43008),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__9581 (
            .O(N__43005),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__9580 (
            .O(N__42998),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__9579 (
            .O(N__42995),
            .I(N__42990));
    CascadeMux I__9578 (
            .O(N__42994),
            .I(N__42987));
    InMux I__9577 (
            .O(N__42993),
            .I(N__42984));
    InMux I__9576 (
            .O(N__42990),
            .I(N__42979));
    InMux I__9575 (
            .O(N__42987),
            .I(N__42979));
    LocalMux I__9574 (
            .O(N__42984),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__9573 (
            .O(N__42979),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__9572 (
            .O(N__42974),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__9571 (
            .O(N__42971),
            .I(N__42966));
    CascadeMux I__9570 (
            .O(N__42970),
            .I(N__42963));
    InMux I__9569 (
            .O(N__42969),
            .I(N__42960));
    InMux I__9568 (
            .O(N__42966),
            .I(N__42955));
    InMux I__9567 (
            .O(N__42963),
            .I(N__42955));
    LocalMux I__9566 (
            .O(N__42960),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__9565 (
            .O(N__42955),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__9564 (
            .O(N__42950),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__9563 (
            .O(N__42947),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__9562 (
            .O(N__42944),
            .I(N__42939));
    InMux I__9561 (
            .O(N__42943),
            .I(N__42934));
    InMux I__9560 (
            .O(N__42942),
            .I(N__42934));
    LocalMux I__9559 (
            .O(N__42939),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__9558 (
            .O(N__42934),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__9557 (
            .O(N__42929),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__9556 (
            .O(N__42926),
            .I(N__42921));
    InMux I__9555 (
            .O(N__42925),
            .I(N__42916));
    InMux I__9554 (
            .O(N__42924),
            .I(N__42916));
    LocalMux I__9553 (
            .O(N__42921),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__9552 (
            .O(N__42916),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__9551 (
            .O(N__42911),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__9550 (
            .O(N__42908),
            .I(N__42903));
    CascadeMux I__9549 (
            .O(N__42907),
            .I(N__42900));
    InMux I__9548 (
            .O(N__42906),
            .I(N__42897));
    InMux I__9547 (
            .O(N__42903),
            .I(N__42892));
    InMux I__9546 (
            .O(N__42900),
            .I(N__42892));
    LocalMux I__9545 (
            .O(N__42897),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__9544 (
            .O(N__42892),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__9543 (
            .O(N__42887),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__9542 (
            .O(N__42884),
            .I(N__42879));
    CascadeMux I__9541 (
            .O(N__42883),
            .I(N__42876));
    InMux I__9540 (
            .O(N__42882),
            .I(N__42873));
    InMux I__9539 (
            .O(N__42879),
            .I(N__42868));
    InMux I__9538 (
            .O(N__42876),
            .I(N__42868));
    LocalMux I__9537 (
            .O(N__42873),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__9536 (
            .O(N__42868),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__9535 (
            .O(N__42863),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__9534 (
            .O(N__42860),
            .I(N__42855));
    InMux I__9533 (
            .O(N__42859),
            .I(N__42852));
    InMux I__9532 (
            .O(N__42858),
            .I(N__42849));
    LocalMux I__9531 (
            .O(N__42855),
            .I(N__42846));
    LocalMux I__9530 (
            .O(N__42852),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__9529 (
            .O(N__42849),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__9528 (
            .O(N__42846),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__9527 (
            .O(N__42839),
            .I(bfn_17_8_0_));
    InMux I__9526 (
            .O(N__42836),
            .I(N__42831));
    InMux I__9525 (
            .O(N__42835),
            .I(N__42828));
    InMux I__9524 (
            .O(N__42834),
            .I(N__42825));
    LocalMux I__9523 (
            .O(N__42831),
            .I(N__42822));
    LocalMux I__9522 (
            .O(N__42828),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__9521 (
            .O(N__42825),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__9520 (
            .O(N__42822),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__9519 (
            .O(N__42815),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__9518 (
            .O(N__42812),
            .I(N__42807));
    CascadeMux I__9517 (
            .O(N__42811),
            .I(N__42804));
    InMux I__9516 (
            .O(N__42810),
            .I(N__42801));
    InMux I__9515 (
            .O(N__42807),
            .I(N__42796));
    InMux I__9514 (
            .O(N__42804),
            .I(N__42796));
    LocalMux I__9513 (
            .O(N__42801),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__9512 (
            .O(N__42796),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__9511 (
            .O(N__42791),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__9510 (
            .O(N__42788),
            .I(N__42783));
    CascadeMux I__9509 (
            .O(N__42787),
            .I(N__42780));
    InMux I__9508 (
            .O(N__42786),
            .I(N__42777));
    InMux I__9507 (
            .O(N__42783),
            .I(N__42772));
    InMux I__9506 (
            .O(N__42780),
            .I(N__42772));
    LocalMux I__9505 (
            .O(N__42777),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__9504 (
            .O(N__42772),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__9503 (
            .O(N__42767),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__9502 (
            .O(N__42764),
            .I(N__42761));
    LocalMux I__9501 (
            .O(N__42761),
            .I(N__42757));
    InMux I__9500 (
            .O(N__42760),
            .I(N__42754));
    Span4Mux_v I__9499 (
            .O(N__42757),
            .I(N__42751));
    LocalMux I__9498 (
            .O(N__42754),
            .I(N__42748));
    Span4Mux_v I__9497 (
            .O(N__42751),
            .I(N__42741));
    Span4Mux_h I__9496 (
            .O(N__42748),
            .I(N__42741));
    InMux I__9495 (
            .O(N__42747),
            .I(N__42738));
    InMux I__9494 (
            .O(N__42746),
            .I(N__42735));
    Odrv4 I__9493 (
            .O(N__42741),
            .I(measured_delay_tr_16));
    LocalMux I__9492 (
            .O(N__42738),
            .I(measured_delay_tr_16));
    LocalMux I__9491 (
            .O(N__42735),
            .I(measured_delay_tr_16));
    CascadeMux I__9490 (
            .O(N__42728),
            .I(N__42725));
    InMux I__9489 (
            .O(N__42725),
            .I(N__42722));
    LocalMux I__9488 (
            .O(N__42722),
            .I(N__42719));
    Span4Mux_v I__9487 (
            .O(N__42719),
            .I(N__42716));
    Span4Mux_h I__9486 (
            .O(N__42716),
            .I(N__42713));
    Odrv4 I__9485 (
            .O(N__42713),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CEMux I__9484 (
            .O(N__42710),
            .I(N__42706));
    CEMux I__9483 (
            .O(N__42709),
            .I(N__42702));
    LocalMux I__9482 (
            .O(N__42706),
            .I(N__42697));
    CEMux I__9481 (
            .O(N__42705),
            .I(N__42694));
    LocalMux I__9480 (
            .O(N__42702),
            .I(N__42691));
    CEMux I__9479 (
            .O(N__42701),
            .I(N__42688));
    CEMux I__9478 (
            .O(N__42700),
            .I(N__42684));
    Span4Mux_v I__9477 (
            .O(N__42697),
            .I(N__42680));
    LocalMux I__9476 (
            .O(N__42694),
            .I(N__42673));
    Span4Mux_v I__9475 (
            .O(N__42691),
            .I(N__42673));
    LocalMux I__9474 (
            .O(N__42688),
            .I(N__42673));
    CEMux I__9473 (
            .O(N__42687),
            .I(N__42670));
    LocalMux I__9472 (
            .O(N__42684),
            .I(N__42667));
    CEMux I__9471 (
            .O(N__42683),
            .I(N__42664));
    Span4Mux_h I__9470 (
            .O(N__42680),
            .I(N__42659));
    Span4Mux_v I__9469 (
            .O(N__42673),
            .I(N__42659));
    LocalMux I__9468 (
            .O(N__42670),
            .I(N__42656));
    Span4Mux_h I__9467 (
            .O(N__42667),
            .I(N__42653));
    LocalMux I__9466 (
            .O(N__42664),
            .I(N__42650));
    Odrv4 I__9465 (
            .O(N__42659),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__9464 (
            .O(N__42656),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__9463 (
            .O(N__42653),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__9462 (
            .O(N__42650),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__9461 (
            .O(N__42641),
            .I(N__42638));
    LocalMux I__9460 (
            .O(N__42638),
            .I(N__42635));
    Span4Mux_h I__9459 (
            .O(N__42635),
            .I(N__42631));
    InMux I__9458 (
            .O(N__42634),
            .I(N__42628));
    Span4Mux_h I__9457 (
            .O(N__42631),
            .I(N__42625));
    LocalMux I__9456 (
            .O(N__42628),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__9455 (
            .O(N__42625),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__9454 (
            .O(N__42620),
            .I(N__42617));
    LocalMux I__9453 (
            .O(N__42617),
            .I(N__42613));
    InMux I__9452 (
            .O(N__42616),
            .I(N__42610));
    Span4Mux_h I__9451 (
            .O(N__42613),
            .I(N__42607));
    LocalMux I__9450 (
            .O(N__42610),
            .I(N__42603));
    Span4Mux_v I__9449 (
            .O(N__42607),
            .I(N__42600));
    InMux I__9448 (
            .O(N__42606),
            .I(N__42597));
    Odrv4 I__9447 (
            .O(N__42603),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__9446 (
            .O(N__42600),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__9445 (
            .O(N__42597),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__9444 (
            .O(N__42590),
            .I(N__42586));
    InMux I__9443 (
            .O(N__42589),
            .I(N__42583));
    LocalMux I__9442 (
            .O(N__42586),
            .I(N__42578));
    LocalMux I__9441 (
            .O(N__42583),
            .I(N__42575));
    InMux I__9440 (
            .O(N__42582),
            .I(N__42572));
    InMux I__9439 (
            .O(N__42581),
            .I(N__42569));
    Span12Mux_h I__9438 (
            .O(N__42578),
            .I(N__42566));
    Span4Mux_v I__9437 (
            .O(N__42575),
            .I(N__42563));
    LocalMux I__9436 (
            .O(N__42572),
            .I(N__42560));
    LocalMux I__9435 (
            .O(N__42569),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__9434 (
            .O(N__42566),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__9433 (
            .O(N__42563),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__9432 (
            .O(N__42560),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__9431 (
            .O(N__42551),
            .I(bfn_17_7_0_));
    InMux I__9430 (
            .O(N__42548),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__9429 (
            .O(N__42545),
            .I(N__42540));
    CascadeMux I__9428 (
            .O(N__42544),
            .I(N__42537));
    InMux I__9427 (
            .O(N__42543),
            .I(N__42534));
    InMux I__9426 (
            .O(N__42540),
            .I(N__42529));
    InMux I__9425 (
            .O(N__42537),
            .I(N__42529));
    LocalMux I__9424 (
            .O(N__42534),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__9423 (
            .O(N__42529),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__9422 (
            .O(N__42524),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    CascadeMux I__9421 (
            .O(N__42521),
            .I(N__42516));
    CascadeMux I__9420 (
            .O(N__42520),
            .I(N__42513));
    InMux I__9419 (
            .O(N__42519),
            .I(N__42510));
    InMux I__9418 (
            .O(N__42516),
            .I(N__42505));
    InMux I__9417 (
            .O(N__42513),
            .I(N__42505));
    LocalMux I__9416 (
            .O(N__42510),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__9415 (
            .O(N__42505),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    CascadeMux I__9414 (
            .O(N__42500),
            .I(N__42496));
    CascadeMux I__9413 (
            .O(N__42499),
            .I(N__42493));
    InMux I__9412 (
            .O(N__42496),
            .I(N__42489));
    InMux I__9411 (
            .O(N__42493),
            .I(N__42484));
    InMux I__9410 (
            .O(N__42492),
            .I(N__42484));
    LocalMux I__9409 (
            .O(N__42489),
            .I(N__42481));
    LocalMux I__9408 (
            .O(N__42484),
            .I(N__42478));
    Span4Mux_h I__9407 (
            .O(N__42481),
            .I(N__42474));
    Span12Mux_v I__9406 (
            .O(N__42478),
            .I(N__42471));
    InMux I__9405 (
            .O(N__42477),
            .I(N__42468));
    Odrv4 I__9404 (
            .O(N__42474),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv12 I__9403 (
            .O(N__42471),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__9402 (
            .O(N__42468),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__9401 (
            .O(N__42461),
            .I(N__42458));
    LocalMux I__9400 (
            .O(N__42458),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    CascadeMux I__9399 (
            .O(N__42455),
            .I(N__42452));
    InMux I__9398 (
            .O(N__42452),
            .I(N__42449));
    LocalMux I__9397 (
            .O(N__42449),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__9396 (
            .O(N__42446),
            .I(N__42443));
    LocalMux I__9395 (
            .O(N__42443),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__9394 (
            .O(N__42440),
            .I(N__42436));
    InMux I__9393 (
            .O(N__42439),
            .I(N__42433));
    LocalMux I__9392 (
            .O(N__42436),
            .I(N__42430));
    LocalMux I__9391 (
            .O(N__42433),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    Odrv12 I__9390 (
            .O(N__42430),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    CascadeMux I__9389 (
            .O(N__42425),
            .I(N__42422));
    InMux I__9388 (
            .O(N__42422),
            .I(N__42419));
    LocalMux I__9387 (
            .O(N__42419),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__9386 (
            .O(N__42416),
            .I(N__42413));
    LocalMux I__9385 (
            .O(N__42413),
            .I(N__42410));
    Odrv4 I__9384 (
            .O(N__42410),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    CascadeMux I__9383 (
            .O(N__42407),
            .I(N__42404));
    InMux I__9382 (
            .O(N__42404),
            .I(N__42401));
    LocalMux I__9381 (
            .O(N__42401),
            .I(N__42398));
    Odrv12 I__9380 (
            .O(N__42398),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__9379 (
            .O(N__42395),
            .I(N__42392));
    LocalMux I__9378 (
            .O(N__42392),
            .I(N__42389));
    Odrv4 I__9377 (
            .O(N__42389),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    InMux I__9376 (
            .O(N__42386),
            .I(N__42383));
    LocalMux I__9375 (
            .O(N__42383),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__9374 (
            .O(N__42380),
            .I(N__42377));
    LocalMux I__9373 (
            .O(N__42377),
            .I(N__42374));
    Odrv12 I__9372 (
            .O(N__42374),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    InMux I__9371 (
            .O(N__42371),
            .I(N__42368));
    LocalMux I__9370 (
            .O(N__42368),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__9369 (
            .O(N__42365),
            .I(N__42362));
    LocalMux I__9368 (
            .O(N__42362),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    CascadeMux I__9367 (
            .O(N__42359),
            .I(N__42356));
    InMux I__9366 (
            .O(N__42356),
            .I(N__42353));
    LocalMux I__9365 (
            .O(N__42353),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    CascadeMux I__9364 (
            .O(N__42350),
            .I(N__42347));
    InMux I__9363 (
            .O(N__42347),
            .I(N__42344));
    LocalMux I__9362 (
            .O(N__42344),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__9361 (
            .O(N__42341),
            .I(N__42338));
    InMux I__9360 (
            .O(N__42338),
            .I(N__42335));
    LocalMux I__9359 (
            .O(N__42335),
            .I(N__42332));
    Odrv4 I__9358 (
            .O(N__42332),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__9357 (
            .O(N__42329),
            .I(N__42326));
    LocalMux I__9356 (
            .O(N__42326),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    InMux I__9355 (
            .O(N__42323),
            .I(N__42320));
    LocalMux I__9354 (
            .O(N__42320),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__9353 (
            .O(N__42317),
            .I(N__42314));
    InMux I__9352 (
            .O(N__42314),
            .I(N__42311));
    LocalMux I__9351 (
            .O(N__42311),
            .I(N__42308));
    Odrv12 I__9350 (
            .O(N__42308),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    CascadeMux I__9349 (
            .O(N__42305),
            .I(N__42302));
    InMux I__9348 (
            .O(N__42302),
            .I(N__42299));
    LocalMux I__9347 (
            .O(N__42299),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    CascadeMux I__9346 (
            .O(N__42296),
            .I(N__42293));
    InMux I__9345 (
            .O(N__42293),
            .I(N__42290));
    LocalMux I__9344 (
            .O(N__42290),
            .I(N__42287));
    Odrv4 I__9343 (
            .O(N__42287),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__9342 (
            .O(N__42284),
            .I(N__42281));
    LocalMux I__9341 (
            .O(N__42281),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    InMux I__9340 (
            .O(N__42278),
            .I(N__42275));
    LocalMux I__9339 (
            .O(N__42275),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__9338 (
            .O(N__42272),
            .I(bfn_16_17_0_));
    InMux I__9337 (
            .O(N__42269),
            .I(N__42266));
    LocalMux I__9336 (
            .O(N__42266),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__9335 (
            .O(N__42263),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__9334 (
            .O(N__42260),
            .I(N__42257));
    LocalMux I__9333 (
            .O(N__42257),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__9332 (
            .O(N__42254),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    CascadeMux I__9331 (
            .O(N__42251),
            .I(N__42248));
    InMux I__9330 (
            .O(N__42248),
            .I(N__42245));
    LocalMux I__9329 (
            .O(N__42245),
            .I(N__42242));
    Span4Mux_v I__9328 (
            .O(N__42242),
            .I(N__42239));
    Odrv4 I__9327 (
            .O(N__42239),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__9326 (
            .O(N__42236),
            .I(N__42233));
    LocalMux I__9325 (
            .O(N__42233),
            .I(N__42230));
    Odrv4 I__9324 (
            .O(N__42230),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__9323 (
            .O(N__42227),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__9322 (
            .O(N__42224),
            .I(N__42221));
    LocalMux I__9321 (
            .O(N__42221),
            .I(N__42218));
    Odrv4 I__9320 (
            .O(N__42218),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__9319 (
            .O(N__42215),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__9318 (
            .O(N__42212),
            .I(N__42209));
    LocalMux I__9317 (
            .O(N__42209),
            .I(N__42206));
    Odrv4 I__9316 (
            .O(N__42206),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__9315 (
            .O(N__42203),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__9314 (
            .O(N__42200),
            .I(N__42197));
    LocalMux I__9313 (
            .O(N__42197),
            .I(N__42194));
    Odrv4 I__9312 (
            .O(N__42194),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__9311 (
            .O(N__42191),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__9310 (
            .O(N__42188),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__9309 (
            .O(N__42185),
            .I(N__42182));
    LocalMux I__9308 (
            .O(N__42182),
            .I(N__42179));
    Odrv4 I__9307 (
            .O(N__42179),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    CascadeMux I__9306 (
            .O(N__42176),
            .I(N__42173));
    InMux I__9305 (
            .O(N__42173),
            .I(N__42170));
    LocalMux I__9304 (
            .O(N__42170),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    InMux I__9303 (
            .O(N__42167),
            .I(N__42164));
    LocalMux I__9302 (
            .O(N__42164),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__9301 (
            .O(N__42161),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__9300 (
            .O(N__42158),
            .I(N__42155));
    LocalMux I__9299 (
            .O(N__42155),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__9298 (
            .O(N__42152),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__9297 (
            .O(N__42149),
            .I(N__42146));
    LocalMux I__9296 (
            .O(N__42146),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__9295 (
            .O(N__42143),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__9294 (
            .O(N__42140),
            .I(N__42137));
    LocalMux I__9293 (
            .O(N__42137),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__9292 (
            .O(N__42134),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    CascadeMux I__9291 (
            .O(N__42131),
            .I(N__42128));
    InMux I__9290 (
            .O(N__42128),
            .I(N__42125));
    LocalMux I__9289 (
            .O(N__42125),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    InMux I__9288 (
            .O(N__42122),
            .I(N__42119));
    LocalMux I__9287 (
            .O(N__42119),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    InMux I__9286 (
            .O(N__42116),
            .I(N__42113));
    LocalMux I__9285 (
            .O(N__42113),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    InMux I__9284 (
            .O(N__42110),
            .I(N__42106));
    InMux I__9283 (
            .O(N__42109),
            .I(N__42103));
    LocalMux I__9282 (
            .O(N__42106),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__9281 (
            .O(N__42103),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__9280 (
            .O(N__42098),
            .I(N__42095));
    LocalMux I__9279 (
            .O(N__42095),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__9278 (
            .O(N__42092),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__9277 (
            .O(N__42089),
            .I(N__42085));
    InMux I__9276 (
            .O(N__42088),
            .I(N__42082));
    LocalMux I__9275 (
            .O(N__42085),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__9274 (
            .O(N__42082),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__9273 (
            .O(N__42077),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__9272 (
            .O(N__42074),
            .I(N__42071));
    LocalMux I__9271 (
            .O(N__42071),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__9270 (
            .O(N__42068),
            .I(N__42065));
    LocalMux I__9269 (
            .O(N__42065),
            .I(N__42061));
    InMux I__9268 (
            .O(N__42064),
            .I(N__42058));
    Span4Mux_h I__9267 (
            .O(N__42061),
            .I(N__42055));
    LocalMux I__9266 (
            .O(N__42058),
            .I(N__42052));
    Span4Mux_v I__9265 (
            .O(N__42055),
            .I(N__42049));
    Odrv12 I__9264 (
            .O(N__42052),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__9263 (
            .O(N__42049),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__9262 (
            .O(N__42044),
            .I(N__42040));
    CascadeMux I__9261 (
            .O(N__42043),
            .I(N__42037));
    InMux I__9260 (
            .O(N__42040),
            .I(N__42034));
    InMux I__9259 (
            .O(N__42037),
            .I(N__42031));
    LocalMux I__9258 (
            .O(N__42034),
            .I(N__42028));
    LocalMux I__9257 (
            .O(N__42031),
            .I(N__42025));
    Span12Mux_s11_h I__9256 (
            .O(N__42028),
            .I(N__42022));
    Span4Mux_v I__9255 (
            .O(N__42025),
            .I(N__42019));
    Odrv12 I__9254 (
            .O(N__42022),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv4 I__9253 (
            .O(N__42019),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__9252 (
            .O(N__42014),
            .I(N__42011));
    LocalMux I__9251 (
            .O(N__42011),
            .I(N__42008));
    Span4Mux_h I__9250 (
            .O(N__42008),
            .I(N__42005));
    Span4Mux_h I__9249 (
            .O(N__42005),
            .I(N__42002));
    Odrv4 I__9248 (
            .O(N__42002),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__9247 (
            .O(N__41999),
            .I(N__41996));
    LocalMux I__9246 (
            .O(N__41996),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    InMux I__9245 (
            .O(N__41993),
            .I(N__41990));
    LocalMux I__9244 (
            .O(N__41990),
            .I(N__41987));
    Span4Mux_h I__9243 (
            .O(N__41987),
            .I(N__41983));
    InMux I__9242 (
            .O(N__41986),
            .I(N__41980));
    Odrv4 I__9241 (
            .O(N__41983),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__9240 (
            .O(N__41980),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__9239 (
            .O(N__41975),
            .I(N__41972));
    LocalMux I__9238 (
            .O(N__41972),
            .I(N__41969));
    Span4Mux_v I__9237 (
            .O(N__41969),
            .I(N__41966));
    Odrv4 I__9236 (
            .O(N__41966),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__9235 (
            .O(N__41963),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__9234 (
            .O(N__41960),
            .I(N__41957));
    LocalMux I__9233 (
            .O(N__41957),
            .I(N__41954));
    Span4Mux_h I__9232 (
            .O(N__41954),
            .I(N__41950));
    InMux I__9231 (
            .O(N__41953),
            .I(N__41947));
    Odrv4 I__9230 (
            .O(N__41950),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__9229 (
            .O(N__41947),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__9228 (
            .O(N__41942),
            .I(N__41939));
    LocalMux I__9227 (
            .O(N__41939),
            .I(N__41936));
    Span4Mux_h I__9226 (
            .O(N__41936),
            .I(N__41933));
    Odrv4 I__9225 (
            .O(N__41933),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__9224 (
            .O(N__41930),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__9223 (
            .O(N__41927),
            .I(N__41924));
    LocalMux I__9222 (
            .O(N__41924),
            .I(N__41921));
    Span4Mux_v I__9221 (
            .O(N__41921),
            .I(N__41917));
    InMux I__9220 (
            .O(N__41920),
            .I(N__41914));
    Odrv4 I__9219 (
            .O(N__41917),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__9218 (
            .O(N__41914),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__9217 (
            .O(N__41909),
            .I(N__41906));
    LocalMux I__9216 (
            .O(N__41906),
            .I(N__41903));
    Span4Mux_h I__9215 (
            .O(N__41903),
            .I(N__41900));
    Odrv4 I__9214 (
            .O(N__41900),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__9213 (
            .O(N__41897),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__9212 (
            .O(N__41894),
            .I(N__41891));
    LocalMux I__9211 (
            .O(N__41891),
            .I(N__41888));
    Span4Mux_v I__9210 (
            .O(N__41888),
            .I(N__41884));
    InMux I__9209 (
            .O(N__41887),
            .I(N__41881));
    Odrv4 I__9208 (
            .O(N__41884),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__9207 (
            .O(N__41881),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__9206 (
            .O(N__41876),
            .I(N__41873));
    LocalMux I__9205 (
            .O(N__41873),
            .I(N__41870));
    Span4Mux_h I__9204 (
            .O(N__41870),
            .I(N__41867));
    Odrv4 I__9203 (
            .O(N__41867),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__9202 (
            .O(N__41864),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__9201 (
            .O(N__41861),
            .I(N__41858));
    LocalMux I__9200 (
            .O(N__41858),
            .I(N__41855));
    Span4Mux_h I__9199 (
            .O(N__41855),
            .I(N__41851));
    InMux I__9198 (
            .O(N__41854),
            .I(N__41848));
    Odrv4 I__9197 (
            .O(N__41851),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__9196 (
            .O(N__41848),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__9195 (
            .O(N__41843),
            .I(N__41840));
    LocalMux I__9194 (
            .O(N__41840),
            .I(N__41837));
    Span4Mux_h I__9193 (
            .O(N__41837),
            .I(N__41834));
    Odrv4 I__9192 (
            .O(N__41834),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__9191 (
            .O(N__41831),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__9190 (
            .O(N__41828),
            .I(N__41825));
    LocalMux I__9189 (
            .O(N__41825),
            .I(N__41822));
    Span4Mux_h I__9188 (
            .O(N__41822),
            .I(N__41818));
    InMux I__9187 (
            .O(N__41821),
            .I(N__41815));
    Odrv4 I__9186 (
            .O(N__41818),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__9185 (
            .O(N__41815),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__9184 (
            .O(N__41810),
            .I(N__41807));
    LocalMux I__9183 (
            .O(N__41807),
            .I(N__41804));
    Span4Mux_h I__9182 (
            .O(N__41804),
            .I(N__41801));
    Odrv4 I__9181 (
            .O(N__41801),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__9180 (
            .O(N__41798),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__9179 (
            .O(N__41795),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__9178 (
            .O(N__41792),
            .I(N__41788));
    InMux I__9177 (
            .O(N__41791),
            .I(N__41785));
    LocalMux I__9176 (
            .O(N__41788),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__9175 (
            .O(N__41785),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__9174 (
            .O(N__41780),
            .I(N__41777));
    LocalMux I__9173 (
            .O(N__41777),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__9172 (
            .O(N__41774),
            .I(bfn_16_13_0_));
    InMux I__9171 (
            .O(N__41771),
            .I(N__41768));
    LocalMux I__9170 (
            .O(N__41768),
            .I(N__41765));
    Odrv4 I__9169 (
            .O(N__41765),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__9168 (
            .O(N__41762),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__9167 (
            .O(N__41759),
            .I(N__41756));
    LocalMux I__9166 (
            .O(N__41756),
            .I(N__41753));
    Span4Mux_h I__9165 (
            .O(N__41753),
            .I(N__41750));
    Odrv4 I__9164 (
            .O(N__41750),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    CascadeMux I__9163 (
            .O(N__41747),
            .I(N__41744));
    InMux I__9162 (
            .O(N__41744),
            .I(N__41740));
    InMux I__9161 (
            .O(N__41743),
            .I(N__41737));
    LocalMux I__9160 (
            .O(N__41740),
            .I(N__41734));
    LocalMux I__9159 (
            .O(N__41737),
            .I(N__41731));
    Odrv4 I__9158 (
            .O(N__41734),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__9157 (
            .O(N__41731),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__9156 (
            .O(N__41726),
            .I(N__41723));
    LocalMux I__9155 (
            .O(N__41723),
            .I(N__41720));
    Odrv4 I__9154 (
            .O(N__41720),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__9153 (
            .O(N__41717),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__9152 (
            .O(N__41714),
            .I(N__41710));
    InMux I__9151 (
            .O(N__41713),
            .I(N__41707));
    LocalMux I__9150 (
            .O(N__41710),
            .I(N__41704));
    LocalMux I__9149 (
            .O(N__41707),
            .I(N__41701));
    Odrv4 I__9148 (
            .O(N__41704),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__9147 (
            .O(N__41701),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__9146 (
            .O(N__41696),
            .I(N__41693));
    LocalMux I__9145 (
            .O(N__41693),
            .I(N__41690));
    Odrv4 I__9144 (
            .O(N__41690),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__9143 (
            .O(N__41687),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__9142 (
            .O(N__41684),
            .I(N__41680));
    InMux I__9141 (
            .O(N__41683),
            .I(N__41677));
    LocalMux I__9140 (
            .O(N__41680),
            .I(N__41674));
    LocalMux I__9139 (
            .O(N__41677),
            .I(N__41671));
    Odrv4 I__9138 (
            .O(N__41674),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv12 I__9137 (
            .O(N__41671),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__9136 (
            .O(N__41666),
            .I(N__41663));
    LocalMux I__9135 (
            .O(N__41663),
            .I(N__41660));
    Odrv4 I__9134 (
            .O(N__41660),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__9133 (
            .O(N__41657),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__9132 (
            .O(N__41654),
            .I(N__41651));
    LocalMux I__9131 (
            .O(N__41651),
            .I(N__41647));
    InMux I__9130 (
            .O(N__41650),
            .I(N__41644));
    Span4Mux_v I__9129 (
            .O(N__41647),
            .I(N__41639));
    LocalMux I__9128 (
            .O(N__41644),
            .I(N__41639));
    Span4Mux_h I__9127 (
            .O(N__41639),
            .I(N__41636));
    Odrv4 I__9126 (
            .O(N__41636),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__9125 (
            .O(N__41633),
            .I(N__41630));
    LocalMux I__9124 (
            .O(N__41630),
            .I(N__41627));
    Odrv4 I__9123 (
            .O(N__41627),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__9122 (
            .O(N__41624),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__9121 (
            .O(N__41621),
            .I(N__41618));
    LocalMux I__9120 (
            .O(N__41618),
            .I(N__41614));
    InMux I__9119 (
            .O(N__41617),
            .I(N__41611));
    Span4Mux_v I__9118 (
            .O(N__41614),
            .I(N__41608));
    LocalMux I__9117 (
            .O(N__41611),
            .I(N__41605));
    Odrv4 I__9116 (
            .O(N__41608),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__9115 (
            .O(N__41605),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__9114 (
            .O(N__41600),
            .I(N__41597));
    LocalMux I__9113 (
            .O(N__41597),
            .I(N__41594));
    Span4Mux_h I__9112 (
            .O(N__41594),
            .I(N__41591));
    Odrv4 I__9111 (
            .O(N__41591),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__9110 (
            .O(N__41588),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__9109 (
            .O(N__41585),
            .I(N__41581));
    InMux I__9108 (
            .O(N__41584),
            .I(N__41578));
    LocalMux I__9107 (
            .O(N__41581),
            .I(N__41575));
    LocalMux I__9106 (
            .O(N__41578),
            .I(N__41572));
    Span4Mux_v I__9105 (
            .O(N__41575),
            .I(N__41569));
    Span4Mux_h I__9104 (
            .O(N__41572),
            .I(N__41566));
    Odrv4 I__9103 (
            .O(N__41569),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__9102 (
            .O(N__41566),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__9101 (
            .O(N__41561),
            .I(N__41558));
    LocalMux I__9100 (
            .O(N__41558),
            .I(N__41555));
    Span4Mux_h I__9099 (
            .O(N__41555),
            .I(N__41552));
    Odrv4 I__9098 (
            .O(N__41552),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__9097 (
            .O(N__41549),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__9096 (
            .O(N__41546),
            .I(N__41543));
    LocalMux I__9095 (
            .O(N__41543),
            .I(N__41539));
    InMux I__9094 (
            .O(N__41542),
            .I(N__41536));
    Odrv4 I__9093 (
            .O(N__41539),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__9092 (
            .O(N__41536),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__9091 (
            .O(N__41531),
            .I(N__41528));
    LocalMux I__9090 (
            .O(N__41528),
            .I(N__41525));
    Odrv4 I__9089 (
            .O(N__41525),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__9088 (
            .O(N__41522),
            .I(bfn_16_12_0_));
    InMux I__9087 (
            .O(N__41519),
            .I(N__41516));
    LocalMux I__9086 (
            .O(N__41516),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__9085 (
            .O(N__41513),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9084 (
            .O(N__41510),
            .I(N__41507));
    LocalMux I__9083 (
            .O(N__41507),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__9082 (
            .O(N__41504),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__9081 (
            .O(N__41501),
            .I(N__41498));
    InMux I__9080 (
            .O(N__41498),
            .I(N__41495));
    LocalMux I__9079 (
            .O(N__41495),
            .I(N__41492));
    Odrv4 I__9078 (
            .O(N__41492),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__9077 (
            .O(N__41489),
            .I(bfn_16_10_0_));
    InMux I__9076 (
            .O(N__41486),
            .I(N__41483));
    LocalMux I__9075 (
            .O(N__41483),
            .I(N__41480));
    Span4Mux_h I__9074 (
            .O(N__41480),
            .I(N__41477));
    Odrv4 I__9073 (
            .O(N__41477),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__9072 (
            .O(N__41474),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__9071 (
            .O(N__41471),
            .I(N__41468));
    LocalMux I__9070 (
            .O(N__41468),
            .I(N__41465));
    Span4Mux_h I__9069 (
            .O(N__41465),
            .I(N__41462));
    Odrv4 I__9068 (
            .O(N__41462),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__9067 (
            .O(N__41459),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__9066 (
            .O(N__41456),
            .I(N__41453));
    InMux I__9065 (
            .O(N__41453),
            .I(N__41450));
    LocalMux I__9064 (
            .O(N__41450),
            .I(N__41447));
    Span4Mux_h I__9063 (
            .O(N__41447),
            .I(N__41444));
    Odrv4 I__9062 (
            .O(N__41444),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__9061 (
            .O(N__41441),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__9060 (
            .O(N__41438),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__9059 (
            .O(N__41435),
            .I(N__41430));
    InMux I__9058 (
            .O(N__41434),
            .I(N__41418));
    InMux I__9057 (
            .O(N__41433),
            .I(N__41418));
    InMux I__9056 (
            .O(N__41430),
            .I(N__41418));
    InMux I__9055 (
            .O(N__41429),
            .I(N__41418));
    CascadeMux I__9054 (
            .O(N__41428),
            .I(N__41414));
    CascadeMux I__9053 (
            .O(N__41427),
            .I(N__41411));
    LocalMux I__9052 (
            .O(N__41418),
            .I(N__41402));
    CascadeMux I__9051 (
            .O(N__41417),
            .I(N__41399));
    InMux I__9050 (
            .O(N__41414),
            .I(N__41396));
    InMux I__9049 (
            .O(N__41411),
            .I(N__41383));
    InMux I__9048 (
            .O(N__41410),
            .I(N__41383));
    InMux I__9047 (
            .O(N__41409),
            .I(N__41383));
    InMux I__9046 (
            .O(N__41408),
            .I(N__41383));
    InMux I__9045 (
            .O(N__41407),
            .I(N__41383));
    InMux I__9044 (
            .O(N__41406),
            .I(N__41383));
    CascadeMux I__9043 (
            .O(N__41405),
            .I(N__41380));
    Span4Mux_v I__9042 (
            .O(N__41402),
            .I(N__41377));
    InMux I__9041 (
            .O(N__41399),
            .I(N__41374));
    LocalMux I__9040 (
            .O(N__41396),
            .I(N__41371));
    LocalMux I__9039 (
            .O(N__41383),
            .I(N__41368));
    InMux I__9038 (
            .O(N__41380),
            .I(N__41365));
    Span4Mux_h I__9037 (
            .O(N__41377),
            .I(N__41360));
    LocalMux I__9036 (
            .O(N__41374),
            .I(N__41360));
    Span4Mux_v I__9035 (
            .O(N__41371),
            .I(N__41353));
    Span4Mux_h I__9034 (
            .O(N__41368),
            .I(N__41353));
    LocalMux I__9033 (
            .O(N__41365),
            .I(N__41353));
    Sp12to4 I__9032 (
            .O(N__41360),
            .I(N__41350));
    Span4Mux_v I__9031 (
            .O(N__41353),
            .I(N__41347));
    Odrv12 I__9030 (
            .O(N__41350),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__9029 (
            .O(N__41347),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    InMux I__9028 (
            .O(N__41342),
            .I(N__41339));
    LocalMux I__9027 (
            .O(N__41339),
            .I(N__41336));
    Span4Mux_h I__9026 (
            .O(N__41336),
            .I(N__41333));
    Odrv4 I__9025 (
            .O(N__41333),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    CascadeMux I__9024 (
            .O(N__41330),
            .I(N__41326));
    InMux I__9023 (
            .O(N__41329),
            .I(N__41323));
    InMux I__9022 (
            .O(N__41326),
            .I(N__41320));
    LocalMux I__9021 (
            .O(N__41323),
            .I(N__41314));
    LocalMux I__9020 (
            .O(N__41320),
            .I(N__41314));
    InMux I__9019 (
            .O(N__41319),
            .I(N__41311));
    Odrv4 I__9018 (
            .O(N__41314),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__9017 (
            .O(N__41311),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__9016 (
            .O(N__41306),
            .I(N__41302));
    InMux I__9015 (
            .O(N__41305),
            .I(N__41299));
    LocalMux I__9014 (
            .O(N__41302),
            .I(N__41296));
    LocalMux I__9013 (
            .O(N__41299),
            .I(N__41293));
    Odrv4 I__9012 (
            .O(N__41296),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__9011 (
            .O(N__41293),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__9010 (
            .O(N__41288),
            .I(N__41285));
    LocalMux I__9009 (
            .O(N__41285),
            .I(N__41282));
    Span4Mux_h I__9008 (
            .O(N__41282),
            .I(N__41277));
    InMux I__9007 (
            .O(N__41281),
            .I(N__41272));
    InMux I__9006 (
            .O(N__41280),
            .I(N__41272));
    Span4Mux_h I__9005 (
            .O(N__41277),
            .I(N__41267));
    LocalMux I__9004 (
            .O(N__41272),
            .I(N__41267));
    Odrv4 I__9003 (
            .O(N__41267),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__9002 (
            .O(N__41264),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__9001 (
            .O(N__41261),
            .I(N__41258));
    LocalMux I__9000 (
            .O(N__41258),
            .I(N__41253));
    InMux I__8999 (
            .O(N__41257),
            .I(N__41248));
    InMux I__8998 (
            .O(N__41256),
            .I(N__41248));
    Span4Mux_v I__8997 (
            .O(N__41253),
            .I(N__41245));
    LocalMux I__8996 (
            .O(N__41248),
            .I(N__41242));
    Odrv4 I__8995 (
            .O(N__41245),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__8994 (
            .O(N__41242),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__8993 (
            .O(N__41237),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__8992 (
            .O(N__41234),
            .I(N__41229));
    CascadeMux I__8991 (
            .O(N__41233),
            .I(N__41226));
    CascadeMux I__8990 (
            .O(N__41232),
            .I(N__41223));
    LocalMux I__8989 (
            .O(N__41229),
            .I(N__41220));
    InMux I__8988 (
            .O(N__41226),
            .I(N__41215));
    InMux I__8987 (
            .O(N__41223),
            .I(N__41215));
    Span12Mux_h I__8986 (
            .O(N__41220),
            .I(N__41212));
    LocalMux I__8985 (
            .O(N__41215),
            .I(N__41209));
    Odrv12 I__8984 (
            .O(N__41212),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    Odrv4 I__8983 (
            .O(N__41209),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__8982 (
            .O(N__41204),
            .I(bfn_16_9_0_));
    InMux I__8981 (
            .O(N__41201),
            .I(N__41198));
    LocalMux I__8980 (
            .O(N__41198),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__8979 (
            .O(N__41195),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__8978 (
            .O(N__41192),
            .I(N__41189));
    LocalMux I__8977 (
            .O(N__41189),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__8976 (
            .O(N__41186),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8975 (
            .O(N__41183),
            .I(N__41180));
    LocalMux I__8974 (
            .O(N__41180),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__8973 (
            .O(N__41177),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__8972 (
            .O(N__41174),
            .I(N__41171));
    InMux I__8971 (
            .O(N__41171),
            .I(N__41168));
    LocalMux I__8970 (
            .O(N__41168),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__8969 (
            .O(N__41165),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8968 (
            .O(N__41162),
            .I(N__41159));
    LocalMux I__8967 (
            .O(N__41159),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__8966 (
            .O(N__41156),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__8965 (
            .O(N__41153),
            .I(N__41150));
    LocalMux I__8964 (
            .O(N__41150),
            .I(N__41146));
    InMux I__8963 (
            .O(N__41149),
            .I(N__41143));
    Span12Mux_v I__8962 (
            .O(N__41146),
            .I(N__41140));
    LocalMux I__8961 (
            .O(N__41143),
            .I(N__41137));
    Odrv12 I__8960 (
            .O(N__41140),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    Odrv12 I__8959 (
            .O(N__41137),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__8958 (
            .O(N__41132),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__8957 (
            .O(N__41129),
            .I(N__41125));
    InMux I__8956 (
            .O(N__41128),
            .I(N__41122));
    LocalMux I__8955 (
            .O(N__41125),
            .I(N__41116));
    LocalMux I__8954 (
            .O(N__41122),
            .I(N__41116));
    InMux I__8953 (
            .O(N__41121),
            .I(N__41113));
    Span4Mux_h I__8952 (
            .O(N__41116),
            .I(N__41108));
    LocalMux I__8951 (
            .O(N__41113),
            .I(N__41105));
    InMux I__8950 (
            .O(N__41112),
            .I(N__41102));
    InMux I__8949 (
            .O(N__41111),
            .I(N__41099));
    Span4Mux_h I__8948 (
            .O(N__41108),
            .I(N__41096));
    Span4Mux_v I__8947 (
            .O(N__41105),
            .I(N__41093));
    LocalMux I__8946 (
            .O(N__41102),
            .I(N__41088));
    LocalMux I__8945 (
            .O(N__41099),
            .I(N__41088));
    Odrv4 I__8944 (
            .O(N__41096),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__8943 (
            .O(N__41093),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv12 I__8942 (
            .O(N__41088),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    InMux I__8941 (
            .O(N__41081),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__8940 (
            .O(N__41078),
            .I(N__41075));
    LocalMux I__8939 (
            .O(N__41075),
            .I(N__41071));
    InMux I__8938 (
            .O(N__41074),
            .I(N__41068));
    Span4Mux_v I__8937 (
            .O(N__41071),
            .I(N__41065));
    LocalMux I__8936 (
            .O(N__41068),
            .I(N__41062));
    Odrv4 I__8935 (
            .O(N__41065),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    Odrv12 I__8934 (
            .O(N__41062),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__8933 (
            .O(N__41057),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__8932 (
            .O(N__41054),
            .I(N__41050));
    InMux I__8931 (
            .O(N__41053),
            .I(N__41047));
    LocalMux I__8930 (
            .O(N__41050),
            .I(N__41042));
    LocalMux I__8929 (
            .O(N__41047),
            .I(N__41042));
    Span12Mux_s7_v I__8928 (
            .O(N__41042),
            .I(N__41039));
    Odrv12 I__8927 (
            .O(N__41039),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__8926 (
            .O(N__41036),
            .I(bfn_16_8_0_));
    InMux I__8925 (
            .O(N__41033),
            .I(N__41029));
    InMux I__8924 (
            .O(N__41032),
            .I(N__41026));
    LocalMux I__8923 (
            .O(N__41029),
            .I(N__41021));
    LocalMux I__8922 (
            .O(N__41026),
            .I(N__41021));
    Span4Mux_v I__8921 (
            .O(N__41021),
            .I(N__41018));
    Span4Mux_h I__8920 (
            .O(N__41018),
            .I(N__41015));
    Odrv4 I__8919 (
            .O(N__41015),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__8918 (
            .O(N__41012),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__8917 (
            .O(N__41009),
            .I(N__41005));
    InMux I__8916 (
            .O(N__41008),
            .I(N__41002));
    InMux I__8915 (
            .O(N__41005),
            .I(N__40999));
    LocalMux I__8914 (
            .O(N__41002),
            .I(N__40994));
    LocalMux I__8913 (
            .O(N__40999),
            .I(N__40994));
    Span4Mux_v I__8912 (
            .O(N__40994),
            .I(N__40991));
    Odrv4 I__8911 (
            .O(N__40991),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__8910 (
            .O(N__40988),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__8909 (
            .O(N__40985),
            .I(N__40980));
    InMux I__8908 (
            .O(N__40984),
            .I(N__40977));
    InMux I__8907 (
            .O(N__40983),
            .I(N__40972));
    LocalMux I__8906 (
            .O(N__40980),
            .I(N__40967));
    LocalMux I__8905 (
            .O(N__40977),
            .I(N__40967));
    InMux I__8904 (
            .O(N__40976),
            .I(N__40964));
    InMux I__8903 (
            .O(N__40975),
            .I(N__40961));
    LocalMux I__8902 (
            .O(N__40972),
            .I(N__40958));
    Span4Mux_v I__8901 (
            .O(N__40967),
            .I(N__40951));
    LocalMux I__8900 (
            .O(N__40964),
            .I(N__40951));
    LocalMux I__8899 (
            .O(N__40961),
            .I(N__40951));
    Span4Mux_v I__8898 (
            .O(N__40958),
            .I(N__40948));
    Span4Mux_h I__8897 (
            .O(N__40951),
            .I(N__40945));
    Odrv4 I__8896 (
            .O(N__40948),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    Odrv4 I__8895 (
            .O(N__40945),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    InMux I__8894 (
            .O(N__40940),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__8893 (
            .O(N__40937),
            .I(N__40929));
    InMux I__8892 (
            .O(N__40936),
            .I(N__40929));
    InMux I__8891 (
            .O(N__40935),
            .I(N__40925));
    CascadeMux I__8890 (
            .O(N__40934),
            .I(N__40921));
    LocalMux I__8889 (
            .O(N__40929),
            .I(N__40918));
    InMux I__8888 (
            .O(N__40928),
            .I(N__40915));
    LocalMux I__8887 (
            .O(N__40925),
            .I(N__40912));
    InMux I__8886 (
            .O(N__40924),
            .I(N__40907));
    InMux I__8885 (
            .O(N__40921),
            .I(N__40907));
    Span4Mux_h I__8884 (
            .O(N__40918),
            .I(N__40904));
    LocalMux I__8883 (
            .O(N__40915),
            .I(N__40901));
    Span4Mux_h I__8882 (
            .O(N__40912),
            .I(N__40896));
    LocalMux I__8881 (
            .O(N__40907),
            .I(N__40896));
    Span4Mux_h I__8880 (
            .O(N__40904),
            .I(N__40893));
    Span4Mux_v I__8879 (
            .O(N__40901),
            .I(N__40888));
    Span4Mux_v I__8878 (
            .O(N__40896),
            .I(N__40888));
    Odrv4 I__8877 (
            .O(N__40893),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv4 I__8876 (
            .O(N__40888),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    InMux I__8875 (
            .O(N__40883),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__8874 (
            .O(N__40880),
            .I(N__40877));
    LocalMux I__8873 (
            .O(N__40877),
            .I(N__40874));
    Span4Mux_v I__8872 (
            .O(N__40874),
            .I(N__40869));
    InMux I__8871 (
            .O(N__40873),
            .I(N__40866));
    InMux I__8870 (
            .O(N__40872),
            .I(N__40863));
    Span4Mux_h I__8869 (
            .O(N__40869),
            .I(N__40856));
    LocalMux I__8868 (
            .O(N__40866),
            .I(N__40856));
    LocalMux I__8867 (
            .O(N__40863),
            .I(N__40856));
    Odrv4 I__8866 (
            .O(N__40856),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__8865 (
            .O(N__40853),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__8864 (
            .O(N__40850),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ));
    InMux I__8863 (
            .O(N__40847),
            .I(N__40844));
    LocalMux I__8862 (
            .O(N__40844),
            .I(N__40841));
    Span4Mux_v I__8861 (
            .O(N__40841),
            .I(N__40838));
    Odrv4 I__8860 (
            .O(N__40838),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ));
    CascadeMux I__8859 (
            .O(N__40835),
            .I(N__40830));
    InMux I__8858 (
            .O(N__40834),
            .I(N__40826));
    InMux I__8857 (
            .O(N__40833),
            .I(N__40823));
    InMux I__8856 (
            .O(N__40830),
            .I(N__40820));
    InMux I__8855 (
            .O(N__40829),
            .I(N__40817));
    LocalMux I__8854 (
            .O(N__40826),
            .I(N__40814));
    LocalMux I__8853 (
            .O(N__40823),
            .I(N__40811));
    LocalMux I__8852 (
            .O(N__40820),
            .I(N__40808));
    LocalMux I__8851 (
            .O(N__40817),
            .I(N__40805));
    Span4Mux_v I__8850 (
            .O(N__40814),
            .I(N__40800));
    Span4Mux_v I__8849 (
            .O(N__40811),
            .I(N__40800));
    Odrv12 I__8848 (
            .O(N__40808),
            .I(\delay_measurement_inst.N_265 ));
    Odrv4 I__8847 (
            .O(N__40805),
            .I(\delay_measurement_inst.N_265 ));
    Odrv4 I__8846 (
            .O(N__40800),
            .I(\delay_measurement_inst.N_265 ));
    InMux I__8845 (
            .O(N__40793),
            .I(N__40790));
    LocalMux I__8844 (
            .O(N__40790),
            .I(N__40787));
    Span4Mux_h I__8843 (
            .O(N__40787),
            .I(N__40783));
    InMux I__8842 (
            .O(N__40786),
            .I(N__40780));
    Odrv4 I__8841 (
            .O(N__40783),
            .I(\delay_measurement_inst.delay_tr_timer.N_287_4 ));
    LocalMux I__8840 (
            .O(N__40780),
            .I(\delay_measurement_inst.delay_tr_timer.N_287_4 ));
    InMux I__8839 (
            .O(N__40775),
            .I(N__40772));
    LocalMux I__8838 (
            .O(N__40772),
            .I(N__40768));
    InMux I__8837 (
            .O(N__40771),
            .I(N__40765));
    Span4Mux_v I__8836 (
            .O(N__40768),
            .I(N__40761));
    LocalMux I__8835 (
            .O(N__40765),
            .I(N__40758));
    InMux I__8834 (
            .O(N__40764),
            .I(N__40755));
    Odrv4 I__8833 (
            .O(N__40761),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    Odrv12 I__8832 (
            .O(N__40758),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    LocalMux I__8831 (
            .O(N__40755),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__8830 (
            .O(N__40748),
            .I(N__40745));
    LocalMux I__8829 (
            .O(N__40745),
            .I(N__40742));
    Span4Mux_v I__8828 (
            .O(N__40742),
            .I(N__40738));
    InMux I__8827 (
            .O(N__40741),
            .I(N__40735));
    Odrv4 I__8826 (
            .O(N__40738),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    LocalMux I__8825 (
            .O(N__40735),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__8824 (
            .O(N__40730),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__8823 (
            .O(N__40727),
            .I(N__40724));
    InMux I__8822 (
            .O(N__40724),
            .I(N__40721));
    LocalMux I__8821 (
            .O(N__40721),
            .I(N__40718));
    Span4Mux_h I__8820 (
            .O(N__40718),
            .I(N__40714));
    InMux I__8819 (
            .O(N__40717),
            .I(N__40711));
    Odrv4 I__8818 (
            .O(N__40714),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    LocalMux I__8817 (
            .O(N__40711),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__8816 (
            .O(N__40706),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__8815 (
            .O(N__40703),
            .I(N__40697));
    CascadeMux I__8814 (
            .O(N__40702),
            .I(N__40693));
    InMux I__8813 (
            .O(N__40701),
            .I(N__40687));
    InMux I__8812 (
            .O(N__40700),
            .I(N__40680));
    InMux I__8811 (
            .O(N__40697),
            .I(N__40680));
    InMux I__8810 (
            .O(N__40696),
            .I(N__40680));
    InMux I__8809 (
            .O(N__40693),
            .I(N__40675));
    InMux I__8808 (
            .O(N__40692),
            .I(N__40675));
    InMux I__8807 (
            .O(N__40691),
            .I(N__40672));
    InMux I__8806 (
            .O(N__40690),
            .I(N__40669));
    LocalMux I__8805 (
            .O(N__40687),
            .I(N__40666));
    LocalMux I__8804 (
            .O(N__40680),
            .I(N__40661));
    LocalMux I__8803 (
            .O(N__40675),
            .I(N__40661));
    LocalMux I__8802 (
            .O(N__40672),
            .I(N__40656));
    LocalMux I__8801 (
            .O(N__40669),
            .I(N__40656));
    Span4Mux_h I__8800 (
            .O(N__40666),
            .I(N__40653));
    Span4Mux_v I__8799 (
            .O(N__40661),
            .I(N__40650));
    Span4Mux_h I__8798 (
            .O(N__40656),
            .I(N__40647));
    Odrv4 I__8797 (
            .O(N__40653),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    Odrv4 I__8796 (
            .O(N__40650),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    Odrv4 I__8795 (
            .O(N__40647),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    InMux I__8794 (
            .O(N__40640),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__8793 (
            .O(N__40637),
            .I(N__40634));
    LocalMux I__8792 (
            .O(N__40634),
            .I(N__40631));
    Span4Mux_v I__8791 (
            .O(N__40631),
            .I(N__40627));
    InMux I__8790 (
            .O(N__40630),
            .I(N__40624));
    Span4Mux_v I__8789 (
            .O(N__40627),
            .I(N__40621));
    LocalMux I__8788 (
            .O(N__40624),
            .I(N__40618));
    Odrv4 I__8787 (
            .O(N__40621),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv12 I__8786 (
            .O(N__40618),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__8785 (
            .O(N__40613),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__8784 (
            .O(N__40610),
            .I(N__40606));
    CascadeMux I__8783 (
            .O(N__40609),
            .I(N__40603));
    InMux I__8782 (
            .O(N__40606),
            .I(N__40598));
    InMux I__8781 (
            .O(N__40603),
            .I(N__40598));
    LocalMux I__8780 (
            .O(N__40598),
            .I(N__40594));
    InMux I__8779 (
            .O(N__40597),
            .I(N__40591));
    Span4Mux_v I__8778 (
            .O(N__40594),
            .I(N__40588));
    LocalMux I__8777 (
            .O(N__40591),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__8776 (
            .O(N__40588),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__8775 (
            .O(N__40583),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__8774 (
            .O(N__40580),
            .I(N__40576));
    CascadeMux I__8773 (
            .O(N__40579),
            .I(N__40573));
    InMux I__8772 (
            .O(N__40576),
            .I(N__40567));
    InMux I__8771 (
            .O(N__40573),
            .I(N__40567));
    InMux I__8770 (
            .O(N__40572),
            .I(N__40564));
    LocalMux I__8769 (
            .O(N__40567),
            .I(N__40561));
    LocalMux I__8768 (
            .O(N__40564),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv12 I__8767 (
            .O(N__40561),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__8766 (
            .O(N__40556),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__8765 (
            .O(N__40553),
            .I(N__40549));
    InMux I__8764 (
            .O(N__40552),
            .I(N__40546));
    LocalMux I__8763 (
            .O(N__40549),
            .I(N__40540));
    LocalMux I__8762 (
            .O(N__40546),
            .I(N__40540));
    InMux I__8761 (
            .O(N__40545),
            .I(N__40537));
    Span4Mux_v I__8760 (
            .O(N__40540),
            .I(N__40534));
    LocalMux I__8759 (
            .O(N__40537),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__8758 (
            .O(N__40534),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__8757 (
            .O(N__40529),
            .I(bfn_15_28_0_));
    InMux I__8756 (
            .O(N__40526),
            .I(N__40522));
    InMux I__8755 (
            .O(N__40525),
            .I(N__40519));
    LocalMux I__8754 (
            .O(N__40522),
            .I(N__40513));
    LocalMux I__8753 (
            .O(N__40519),
            .I(N__40513));
    InMux I__8752 (
            .O(N__40518),
            .I(N__40510));
    Span4Mux_v I__8751 (
            .O(N__40513),
            .I(N__40507));
    LocalMux I__8750 (
            .O(N__40510),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__8749 (
            .O(N__40507),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__8748 (
            .O(N__40502),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__8747 (
            .O(N__40499),
            .I(N__40495));
    CascadeMux I__8746 (
            .O(N__40498),
            .I(N__40492));
    InMux I__8745 (
            .O(N__40495),
            .I(N__40487));
    InMux I__8744 (
            .O(N__40492),
            .I(N__40487));
    LocalMux I__8743 (
            .O(N__40487),
            .I(N__40483));
    InMux I__8742 (
            .O(N__40486),
            .I(N__40480));
    Span4Mux_h I__8741 (
            .O(N__40483),
            .I(N__40477));
    LocalMux I__8740 (
            .O(N__40480),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__8739 (
            .O(N__40477),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__8738 (
            .O(N__40472),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__8737 (
            .O(N__40469),
            .I(N__40465));
    CascadeMux I__8736 (
            .O(N__40468),
            .I(N__40462));
    InMux I__8735 (
            .O(N__40465),
            .I(N__40457));
    InMux I__8734 (
            .O(N__40462),
            .I(N__40457));
    LocalMux I__8733 (
            .O(N__40457),
            .I(N__40453));
    InMux I__8732 (
            .O(N__40456),
            .I(N__40450));
    Span4Mux_h I__8731 (
            .O(N__40453),
            .I(N__40447));
    LocalMux I__8730 (
            .O(N__40450),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__8729 (
            .O(N__40447),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__8728 (
            .O(N__40442),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__8727 (
            .O(N__40439),
            .I(N__40436));
    LocalMux I__8726 (
            .O(N__40436),
            .I(N__40432));
    InMux I__8725 (
            .O(N__40435),
            .I(N__40429));
    Span4Mux_h I__8724 (
            .O(N__40432),
            .I(N__40426));
    LocalMux I__8723 (
            .O(N__40429),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__8722 (
            .O(N__40426),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__8721 (
            .O(N__40421),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__8720 (
            .O(N__40418),
            .I(N__40396));
    InMux I__8719 (
            .O(N__40417),
            .I(N__40396));
    InMux I__8718 (
            .O(N__40416),
            .I(N__40387));
    InMux I__8717 (
            .O(N__40415),
            .I(N__40387));
    InMux I__8716 (
            .O(N__40414),
            .I(N__40387));
    InMux I__8715 (
            .O(N__40413),
            .I(N__40387));
    InMux I__8714 (
            .O(N__40412),
            .I(N__40366));
    InMux I__8713 (
            .O(N__40411),
            .I(N__40366));
    InMux I__8712 (
            .O(N__40410),
            .I(N__40366));
    InMux I__8711 (
            .O(N__40409),
            .I(N__40366));
    InMux I__8710 (
            .O(N__40408),
            .I(N__40357));
    InMux I__8709 (
            .O(N__40407),
            .I(N__40357));
    InMux I__8708 (
            .O(N__40406),
            .I(N__40357));
    InMux I__8707 (
            .O(N__40405),
            .I(N__40357));
    InMux I__8706 (
            .O(N__40404),
            .I(N__40348));
    InMux I__8705 (
            .O(N__40403),
            .I(N__40348));
    InMux I__8704 (
            .O(N__40402),
            .I(N__40348));
    InMux I__8703 (
            .O(N__40401),
            .I(N__40348));
    LocalMux I__8702 (
            .O(N__40396),
            .I(N__40343));
    LocalMux I__8701 (
            .O(N__40387),
            .I(N__40343));
    InMux I__8700 (
            .O(N__40386),
            .I(N__40334));
    InMux I__8699 (
            .O(N__40385),
            .I(N__40334));
    InMux I__8698 (
            .O(N__40384),
            .I(N__40334));
    InMux I__8697 (
            .O(N__40383),
            .I(N__40334));
    InMux I__8696 (
            .O(N__40382),
            .I(N__40325));
    InMux I__8695 (
            .O(N__40381),
            .I(N__40325));
    InMux I__8694 (
            .O(N__40380),
            .I(N__40325));
    InMux I__8693 (
            .O(N__40379),
            .I(N__40325));
    InMux I__8692 (
            .O(N__40378),
            .I(N__40316));
    InMux I__8691 (
            .O(N__40377),
            .I(N__40316));
    InMux I__8690 (
            .O(N__40376),
            .I(N__40316));
    InMux I__8689 (
            .O(N__40375),
            .I(N__40316));
    LocalMux I__8688 (
            .O(N__40366),
            .I(N__40307));
    LocalMux I__8687 (
            .O(N__40357),
            .I(N__40307));
    LocalMux I__8686 (
            .O(N__40348),
            .I(N__40307));
    Span4Mux_s3_v I__8685 (
            .O(N__40343),
            .I(N__40307));
    LocalMux I__8684 (
            .O(N__40334),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__8683 (
            .O(N__40325),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__8682 (
            .O(N__40316),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__8681 (
            .O(N__40307),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__8680 (
            .O(N__40298),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__8679 (
            .O(N__40295),
            .I(N__40292));
    LocalMux I__8678 (
            .O(N__40292),
            .I(N__40288));
    InMux I__8677 (
            .O(N__40291),
            .I(N__40285));
    Span4Mux_h I__8676 (
            .O(N__40288),
            .I(N__40282));
    LocalMux I__8675 (
            .O(N__40285),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__8674 (
            .O(N__40282),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__8673 (
            .O(N__40277),
            .I(N__40265));
    CEMux I__8672 (
            .O(N__40276),
            .I(N__40265));
    CEMux I__8671 (
            .O(N__40275),
            .I(N__40265));
    CEMux I__8670 (
            .O(N__40274),
            .I(N__40265));
    GlobalMux I__8669 (
            .O(N__40265),
            .I(N__40262));
    gio2CtrlBuf I__8668 (
            .O(N__40262),
            .I(\current_shift_inst.timer_s1.N_181_i_g ));
    CascadeMux I__8667 (
            .O(N__40259),
            .I(N__40255));
    CascadeMux I__8666 (
            .O(N__40258),
            .I(N__40252));
    InMux I__8665 (
            .O(N__40255),
            .I(N__40246));
    InMux I__8664 (
            .O(N__40252),
            .I(N__40246));
    InMux I__8663 (
            .O(N__40251),
            .I(N__40243));
    LocalMux I__8662 (
            .O(N__40246),
            .I(N__40240));
    LocalMux I__8661 (
            .O(N__40243),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv12 I__8660 (
            .O(N__40240),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__8659 (
            .O(N__40235),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__8658 (
            .O(N__40232),
            .I(N__40228));
    CascadeMux I__8657 (
            .O(N__40231),
            .I(N__40225));
    InMux I__8656 (
            .O(N__40228),
            .I(N__40220));
    InMux I__8655 (
            .O(N__40225),
            .I(N__40220));
    LocalMux I__8654 (
            .O(N__40220),
            .I(N__40216));
    InMux I__8653 (
            .O(N__40219),
            .I(N__40213));
    Span4Mux_v I__8652 (
            .O(N__40216),
            .I(N__40210));
    LocalMux I__8651 (
            .O(N__40213),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__8650 (
            .O(N__40210),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__8649 (
            .O(N__40205),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__8648 (
            .O(N__40202),
            .I(N__40198));
    InMux I__8647 (
            .O(N__40201),
            .I(N__40195));
    LocalMux I__8646 (
            .O(N__40198),
            .I(N__40189));
    LocalMux I__8645 (
            .O(N__40195),
            .I(N__40189));
    InMux I__8644 (
            .O(N__40194),
            .I(N__40186));
    Span4Mux_v I__8643 (
            .O(N__40189),
            .I(N__40183));
    LocalMux I__8642 (
            .O(N__40186),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__8641 (
            .O(N__40183),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__8640 (
            .O(N__40178),
            .I(bfn_15_27_0_));
    InMux I__8639 (
            .O(N__40175),
            .I(N__40171));
    InMux I__8638 (
            .O(N__40174),
            .I(N__40168));
    LocalMux I__8637 (
            .O(N__40171),
            .I(N__40164));
    LocalMux I__8636 (
            .O(N__40168),
            .I(N__40161));
    InMux I__8635 (
            .O(N__40167),
            .I(N__40158));
    Span4Mux_v I__8634 (
            .O(N__40164),
            .I(N__40153));
    Span4Mux_v I__8633 (
            .O(N__40161),
            .I(N__40153));
    LocalMux I__8632 (
            .O(N__40158),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__8631 (
            .O(N__40153),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__8630 (
            .O(N__40148),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__8629 (
            .O(N__40145),
            .I(N__40141));
    CascadeMux I__8628 (
            .O(N__40144),
            .I(N__40138));
    InMux I__8627 (
            .O(N__40141),
            .I(N__40133));
    InMux I__8626 (
            .O(N__40138),
            .I(N__40133));
    LocalMux I__8625 (
            .O(N__40133),
            .I(N__40129));
    InMux I__8624 (
            .O(N__40132),
            .I(N__40126));
    Span4Mux_h I__8623 (
            .O(N__40129),
            .I(N__40123));
    LocalMux I__8622 (
            .O(N__40126),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__8621 (
            .O(N__40123),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__8620 (
            .O(N__40118),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__8619 (
            .O(N__40115),
            .I(N__40111));
    CascadeMux I__8618 (
            .O(N__40114),
            .I(N__40108));
    InMux I__8617 (
            .O(N__40111),
            .I(N__40103));
    InMux I__8616 (
            .O(N__40108),
            .I(N__40103));
    LocalMux I__8615 (
            .O(N__40103),
            .I(N__40099));
    InMux I__8614 (
            .O(N__40102),
            .I(N__40096));
    Span4Mux_h I__8613 (
            .O(N__40099),
            .I(N__40093));
    LocalMux I__8612 (
            .O(N__40096),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__8611 (
            .O(N__40093),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__8610 (
            .O(N__40088),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__8609 (
            .O(N__40085),
            .I(N__40078));
    InMux I__8608 (
            .O(N__40084),
            .I(N__40078));
    InMux I__8607 (
            .O(N__40083),
            .I(N__40075));
    LocalMux I__8606 (
            .O(N__40078),
            .I(N__40072));
    LocalMux I__8605 (
            .O(N__40075),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv12 I__8604 (
            .O(N__40072),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__8603 (
            .O(N__40067),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__8602 (
            .O(N__40064),
            .I(N__40058));
    InMux I__8601 (
            .O(N__40063),
            .I(N__40058));
    LocalMux I__8600 (
            .O(N__40058),
            .I(N__40054));
    InMux I__8599 (
            .O(N__40057),
            .I(N__40051));
    Span4Mux_h I__8598 (
            .O(N__40054),
            .I(N__40048));
    LocalMux I__8597 (
            .O(N__40051),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__8596 (
            .O(N__40048),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__8595 (
            .O(N__40043),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__8594 (
            .O(N__40040),
            .I(N__40034));
    InMux I__8593 (
            .O(N__40039),
            .I(N__40034));
    LocalMux I__8592 (
            .O(N__40034),
            .I(N__40030));
    InMux I__8591 (
            .O(N__40033),
            .I(N__40027));
    Span4Mux_v I__8590 (
            .O(N__40030),
            .I(N__40024));
    LocalMux I__8589 (
            .O(N__40027),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__8588 (
            .O(N__40024),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__8587 (
            .O(N__40019),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__8586 (
            .O(N__40016),
            .I(N__40010));
    InMux I__8585 (
            .O(N__40015),
            .I(N__40010));
    LocalMux I__8584 (
            .O(N__40010),
            .I(N__40006));
    InMux I__8583 (
            .O(N__40009),
            .I(N__40003));
    Span4Mux_v I__8582 (
            .O(N__40006),
            .I(N__40000));
    LocalMux I__8581 (
            .O(N__40003),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__8580 (
            .O(N__40000),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__8579 (
            .O(N__39995),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__8578 (
            .O(N__39992),
            .I(N__39988));
    InMux I__8577 (
            .O(N__39991),
            .I(N__39985));
    InMux I__8576 (
            .O(N__39988),
            .I(N__39982));
    LocalMux I__8575 (
            .O(N__39985),
            .I(N__39976));
    LocalMux I__8574 (
            .O(N__39982),
            .I(N__39976));
    InMux I__8573 (
            .O(N__39981),
            .I(N__39973));
    Span4Mux_v I__8572 (
            .O(N__39976),
            .I(N__39970));
    LocalMux I__8571 (
            .O(N__39973),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__8570 (
            .O(N__39970),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__8569 (
            .O(N__39965),
            .I(bfn_15_26_0_));
    CascadeMux I__8568 (
            .O(N__39962),
            .I(N__39958));
    InMux I__8567 (
            .O(N__39961),
            .I(N__39955));
    InMux I__8566 (
            .O(N__39958),
            .I(N__39952));
    LocalMux I__8565 (
            .O(N__39955),
            .I(N__39946));
    LocalMux I__8564 (
            .O(N__39952),
            .I(N__39946));
    InMux I__8563 (
            .O(N__39951),
            .I(N__39943));
    Span4Mux_v I__8562 (
            .O(N__39946),
            .I(N__39940));
    LocalMux I__8561 (
            .O(N__39943),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__8560 (
            .O(N__39940),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__8559 (
            .O(N__39935),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__8558 (
            .O(N__39932),
            .I(N__39928));
    CascadeMux I__8557 (
            .O(N__39931),
            .I(N__39925));
    InMux I__8556 (
            .O(N__39928),
            .I(N__39920));
    InMux I__8555 (
            .O(N__39925),
            .I(N__39920));
    LocalMux I__8554 (
            .O(N__39920),
            .I(N__39916));
    InMux I__8553 (
            .O(N__39919),
            .I(N__39913));
    Span4Mux_h I__8552 (
            .O(N__39916),
            .I(N__39910));
    LocalMux I__8551 (
            .O(N__39913),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__8550 (
            .O(N__39910),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__8549 (
            .O(N__39905),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__8548 (
            .O(N__39902),
            .I(N__39898));
    CascadeMux I__8547 (
            .O(N__39901),
            .I(N__39895));
    InMux I__8546 (
            .O(N__39898),
            .I(N__39889));
    InMux I__8545 (
            .O(N__39895),
            .I(N__39889));
    InMux I__8544 (
            .O(N__39894),
            .I(N__39886));
    LocalMux I__8543 (
            .O(N__39889),
            .I(N__39883));
    LocalMux I__8542 (
            .O(N__39886),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv12 I__8541 (
            .O(N__39883),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__8540 (
            .O(N__39878),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__8539 (
            .O(N__39875),
            .I(N__39868));
    InMux I__8538 (
            .O(N__39874),
            .I(N__39868));
    InMux I__8537 (
            .O(N__39873),
            .I(N__39865));
    LocalMux I__8536 (
            .O(N__39868),
            .I(N__39862));
    LocalMux I__8535 (
            .O(N__39865),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv12 I__8534 (
            .O(N__39862),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__8533 (
            .O(N__39857),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__8532 (
            .O(N__39854),
            .I(N__39847));
    InMux I__8531 (
            .O(N__39853),
            .I(N__39847));
    InMux I__8530 (
            .O(N__39852),
            .I(N__39844));
    LocalMux I__8529 (
            .O(N__39847),
            .I(N__39841));
    LocalMux I__8528 (
            .O(N__39844),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv12 I__8527 (
            .O(N__39841),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__8526 (
            .O(N__39836),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__8525 (
            .O(N__39833),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__8524 (
            .O(N__39830),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__8523 (
            .O(N__39827),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__8522 (
            .O(N__39824),
            .I(bfn_15_25_0_));
    InMux I__8521 (
            .O(N__39821),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__8520 (
            .O(N__39818),
            .I(N__39811));
    InMux I__8519 (
            .O(N__39817),
            .I(N__39811));
    InMux I__8518 (
            .O(N__39816),
            .I(N__39808));
    LocalMux I__8517 (
            .O(N__39811),
            .I(N__39805));
    LocalMux I__8516 (
            .O(N__39808),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__8515 (
            .O(N__39805),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__8514 (
            .O(N__39800),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__8513 (
            .O(N__39797),
            .I(N__39791));
    InMux I__8512 (
            .O(N__39796),
            .I(N__39791));
    LocalMux I__8511 (
            .O(N__39791),
            .I(N__39787));
    InMux I__8510 (
            .O(N__39790),
            .I(N__39784));
    Span4Mux_h I__8509 (
            .O(N__39787),
            .I(N__39781));
    LocalMux I__8508 (
            .O(N__39784),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__8507 (
            .O(N__39781),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__8506 (
            .O(N__39776),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__8505 (
            .O(N__39773),
            .I(N__39769));
    CascadeMux I__8504 (
            .O(N__39772),
            .I(N__39766));
    InMux I__8503 (
            .O(N__39769),
            .I(N__39760));
    InMux I__8502 (
            .O(N__39766),
            .I(N__39760));
    InMux I__8501 (
            .O(N__39765),
            .I(N__39757));
    LocalMux I__8500 (
            .O(N__39760),
            .I(N__39754));
    LocalMux I__8499 (
            .O(N__39757),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv12 I__8498 (
            .O(N__39754),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__8497 (
            .O(N__39749),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__8496 (
            .O(N__39746),
            .I(N__39742));
    CascadeMux I__8495 (
            .O(N__39745),
            .I(N__39739));
    InMux I__8494 (
            .O(N__39742),
            .I(N__39733));
    InMux I__8493 (
            .O(N__39739),
            .I(N__39733));
    InMux I__8492 (
            .O(N__39738),
            .I(N__39730));
    LocalMux I__8491 (
            .O(N__39733),
            .I(N__39727));
    LocalMux I__8490 (
            .O(N__39730),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv12 I__8489 (
            .O(N__39727),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__8488 (
            .O(N__39722),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__8487 (
            .O(N__39719),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__8486 (
            .O(N__39716),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__8485 (
            .O(N__39713),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__8484 (
            .O(N__39710),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__8483 (
            .O(N__39707),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__8482 (
            .O(N__39704),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__8481 (
            .O(N__39701),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__8480 (
            .O(N__39698),
            .I(bfn_15_24_0_));
    InMux I__8479 (
            .O(N__39695),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__8478 (
            .O(N__39692),
            .I(bfn_15_22_0_));
    InMux I__8477 (
            .O(N__39689),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__8476 (
            .O(N__39686),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__8475 (
            .O(N__39683),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__8474 (
            .O(N__39680),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__8473 (
            .O(N__39677),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__8472 (
            .O(N__39674),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__8471 (
            .O(N__39671),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__8470 (
            .O(N__39668),
            .I(bfn_15_23_0_));
    InMux I__8469 (
            .O(N__39665),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__8468 (
            .O(N__39662),
            .I(N__39659));
    LocalMux I__8467 (
            .O(N__39659),
            .I(N__39656));
    Span4Mux_h I__8466 (
            .O(N__39656),
            .I(N__39653));
    Odrv4 I__8465 (
            .O(N__39653),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__8464 (
            .O(N__39650),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__8463 (
            .O(N__39647),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__8462 (
            .O(N__39644),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__8461 (
            .O(N__39641),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__8460 (
            .O(N__39638),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__8459 (
            .O(N__39635),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__8458 (
            .O(N__39632),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__8457 (
            .O(N__39629),
            .I(N__39626));
    InMux I__8456 (
            .O(N__39626),
            .I(N__39623));
    LocalMux I__8455 (
            .O(N__39623),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__8454 (
            .O(N__39620),
            .I(N__39617));
    LocalMux I__8453 (
            .O(N__39617),
            .I(N__39614));
    Span4Mux_v I__8452 (
            .O(N__39614),
            .I(N__39611));
    Odrv4 I__8451 (
            .O(N__39611),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__8450 (
            .O(N__39608),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__8449 (
            .O(N__39605),
            .I(N__39602));
    LocalMux I__8448 (
            .O(N__39602),
            .I(N__39599));
    Span4Mux_h I__8447 (
            .O(N__39599),
            .I(N__39596));
    Odrv4 I__8446 (
            .O(N__39596),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__8445 (
            .O(N__39593),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    CascadeMux I__8444 (
            .O(N__39590),
            .I(N__39587));
    InMux I__8443 (
            .O(N__39587),
            .I(N__39584));
    LocalMux I__8442 (
            .O(N__39584),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__8441 (
            .O(N__39581),
            .I(N__39578));
    LocalMux I__8440 (
            .O(N__39578),
            .I(N__39575));
    Span4Mux_h I__8439 (
            .O(N__39575),
            .I(N__39572));
    Odrv4 I__8438 (
            .O(N__39572),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__8437 (
            .O(N__39569),
            .I(bfn_15_20_0_));
    InMux I__8436 (
            .O(N__39566),
            .I(N__39563));
    LocalMux I__8435 (
            .O(N__39563),
            .I(N__39560));
    Span4Mux_h I__8434 (
            .O(N__39560),
            .I(N__39557));
    Odrv4 I__8433 (
            .O(N__39557),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__8432 (
            .O(N__39554),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__8431 (
            .O(N__39551),
            .I(N__39548));
    LocalMux I__8430 (
            .O(N__39548),
            .I(N__39545));
    Span4Mux_h I__8429 (
            .O(N__39545),
            .I(N__39542));
    Odrv4 I__8428 (
            .O(N__39542),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__8427 (
            .O(N__39539),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__8426 (
            .O(N__39536),
            .I(N__39533));
    LocalMux I__8425 (
            .O(N__39533),
            .I(N__39530));
    Span4Mux_v I__8424 (
            .O(N__39530),
            .I(N__39527));
    Odrv4 I__8423 (
            .O(N__39527),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__8422 (
            .O(N__39524),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__8421 (
            .O(N__39521),
            .I(N__39518));
    LocalMux I__8420 (
            .O(N__39518),
            .I(N__39515));
    Odrv4 I__8419 (
            .O(N__39515),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__8418 (
            .O(N__39512),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__8417 (
            .O(N__39509),
            .I(N__39506));
    LocalMux I__8416 (
            .O(N__39506),
            .I(N__39503));
    Odrv12 I__8415 (
            .O(N__39503),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__8414 (
            .O(N__39500),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__8413 (
            .O(N__39497),
            .I(N__39494));
    LocalMux I__8412 (
            .O(N__39494),
            .I(N__39491));
    Odrv12 I__8411 (
            .O(N__39491),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__8410 (
            .O(N__39488),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__8409 (
            .O(N__39485),
            .I(N__39482));
    LocalMux I__8408 (
            .O(N__39482),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    InMux I__8407 (
            .O(N__39479),
            .I(N__39476));
    LocalMux I__8406 (
            .O(N__39476),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    CascadeMux I__8405 (
            .O(N__39473),
            .I(N__39470));
    InMux I__8404 (
            .O(N__39470),
            .I(N__39467));
    LocalMux I__8403 (
            .O(N__39467),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    InMux I__8402 (
            .O(N__39464),
            .I(N__39461));
    LocalMux I__8401 (
            .O(N__39461),
            .I(N__39458));
    Odrv4 I__8400 (
            .O(N__39458),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__8399 (
            .O(N__39455),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__8398 (
            .O(N__39452),
            .I(N__39449));
    LocalMux I__8397 (
            .O(N__39449),
            .I(N__39446));
    Odrv12 I__8396 (
            .O(N__39446),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__8395 (
            .O(N__39443),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__8394 (
            .O(N__39440),
            .I(N__39437));
    LocalMux I__8393 (
            .O(N__39437),
            .I(N__39434));
    Span4Mux_v I__8392 (
            .O(N__39434),
            .I(N__39431));
    Odrv4 I__8391 (
            .O(N__39431),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    InMux I__8390 (
            .O(N__39428),
            .I(N__39425));
    LocalMux I__8389 (
            .O(N__39425),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    InMux I__8388 (
            .O(N__39422),
            .I(N__39419));
    LocalMux I__8387 (
            .O(N__39419),
            .I(N__39416));
    Odrv12 I__8386 (
            .O(N__39416),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    InMux I__8385 (
            .O(N__39413),
            .I(N__39410));
    LocalMux I__8384 (
            .O(N__39410),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    InMux I__8383 (
            .O(N__39407),
            .I(N__39404));
    LocalMux I__8382 (
            .O(N__39404),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__8381 (
            .O(N__39401),
            .I(N__39398));
    LocalMux I__8380 (
            .O(N__39398),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__8379 (
            .O(N__39395),
            .I(N__39392));
    LocalMux I__8378 (
            .O(N__39392),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__8377 (
            .O(N__39389),
            .I(N__39386));
    LocalMux I__8376 (
            .O(N__39386),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__8375 (
            .O(N__39383),
            .I(N__39380));
    LocalMux I__8374 (
            .O(N__39380),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__8373 (
            .O(N__39377),
            .I(N__39374));
    LocalMux I__8372 (
            .O(N__39374),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__8371 (
            .O(N__39371),
            .I(N__39368));
    InMux I__8370 (
            .O(N__39368),
            .I(N__39365));
    LocalMux I__8369 (
            .O(N__39365),
            .I(N__39362));
    Odrv4 I__8368 (
            .O(N__39362),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    InMux I__8367 (
            .O(N__39359),
            .I(N__39356));
    LocalMux I__8366 (
            .O(N__39356),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__8365 (
            .O(N__39353),
            .I(N__39350));
    LocalMux I__8364 (
            .O(N__39350),
            .I(N__39347));
    Odrv4 I__8363 (
            .O(N__39347),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    CascadeMux I__8362 (
            .O(N__39344),
            .I(N__39341));
    InMux I__8361 (
            .O(N__39341),
            .I(N__39338));
    LocalMux I__8360 (
            .O(N__39338),
            .I(N__39335));
    Odrv4 I__8359 (
            .O(N__39335),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__8358 (
            .O(N__39332),
            .I(N__39328));
    InMux I__8357 (
            .O(N__39331),
            .I(N__39323));
    LocalMux I__8356 (
            .O(N__39328),
            .I(N__39320));
    InMux I__8355 (
            .O(N__39327),
            .I(N__39317));
    CascadeMux I__8354 (
            .O(N__39326),
            .I(N__39314));
    LocalMux I__8353 (
            .O(N__39323),
            .I(N__39311));
    Span4Mux_h I__8352 (
            .O(N__39320),
            .I(N__39308));
    LocalMux I__8351 (
            .O(N__39317),
            .I(N__39305));
    InMux I__8350 (
            .O(N__39314),
            .I(N__39302));
    Span4Mux_v I__8349 (
            .O(N__39311),
            .I(N__39297));
    Span4Mux_v I__8348 (
            .O(N__39308),
            .I(N__39297));
    Span12Mux_v I__8347 (
            .O(N__39305),
            .I(N__39294));
    LocalMux I__8346 (
            .O(N__39302),
            .I(measured_delay_tr_7));
    Odrv4 I__8345 (
            .O(N__39297),
            .I(measured_delay_tr_7));
    Odrv12 I__8344 (
            .O(N__39294),
            .I(measured_delay_tr_7));
    InMux I__8343 (
            .O(N__39287),
            .I(N__39281));
    InMux I__8342 (
            .O(N__39286),
            .I(N__39281));
    LocalMux I__8341 (
            .O(N__39281),
            .I(N__39278));
    Span4Mux_v I__8340 (
            .O(N__39278),
            .I(N__39274));
    InMux I__8339 (
            .O(N__39277),
            .I(N__39271));
    Span4Mux_v I__8338 (
            .O(N__39274),
            .I(N__39268));
    LocalMux I__8337 (
            .O(N__39271),
            .I(N__39265));
    Odrv4 I__8336 (
            .O(N__39268),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    Odrv4 I__8335 (
            .O(N__39265),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    CascadeMux I__8334 (
            .O(N__39260),
            .I(N__39256));
    CascadeMux I__8333 (
            .O(N__39259),
            .I(N__39253));
    InMux I__8332 (
            .O(N__39256),
            .I(N__39244));
    InMux I__8331 (
            .O(N__39253),
            .I(N__39237));
    InMux I__8330 (
            .O(N__39252),
            .I(N__39237));
    InMux I__8329 (
            .O(N__39251),
            .I(N__39237));
    InMux I__8328 (
            .O(N__39250),
            .I(N__39232));
    InMux I__8327 (
            .O(N__39249),
            .I(N__39232));
    InMux I__8326 (
            .O(N__39248),
            .I(N__39227));
    InMux I__8325 (
            .O(N__39247),
            .I(N__39227));
    LocalMux I__8324 (
            .O(N__39244),
            .I(N__39220));
    LocalMux I__8323 (
            .O(N__39237),
            .I(N__39220));
    LocalMux I__8322 (
            .O(N__39232),
            .I(N__39220));
    LocalMux I__8321 (
            .O(N__39227),
            .I(N__39217));
    Span4Mux_v I__8320 (
            .O(N__39220),
            .I(N__39214));
    Span12Mux_v I__8319 (
            .O(N__39217),
            .I(N__39211));
    Odrv4 I__8318 (
            .O(N__39214),
            .I(\delay_measurement_inst.N_267 ));
    Odrv12 I__8317 (
            .O(N__39211),
            .I(\delay_measurement_inst.N_267 ));
    InMux I__8316 (
            .O(N__39206),
            .I(N__39201));
    InMux I__8315 (
            .O(N__39205),
            .I(N__39198));
    InMux I__8314 (
            .O(N__39204),
            .I(N__39195));
    LocalMux I__8313 (
            .O(N__39201),
            .I(N__39190));
    LocalMux I__8312 (
            .O(N__39198),
            .I(N__39190));
    LocalMux I__8311 (
            .O(N__39195),
            .I(N__39184));
    Span4Mux_h I__8310 (
            .O(N__39190),
            .I(N__39184));
    CascadeMux I__8309 (
            .O(N__39189),
            .I(N__39181));
    Span4Mux_v I__8308 (
            .O(N__39184),
            .I(N__39178));
    InMux I__8307 (
            .O(N__39181),
            .I(N__39175));
    Span4Mux_v I__8306 (
            .O(N__39178),
            .I(N__39172));
    LocalMux I__8305 (
            .O(N__39175),
            .I(measured_delay_tr_8));
    Odrv4 I__8304 (
            .O(N__39172),
            .I(measured_delay_tr_8));
    InMux I__8303 (
            .O(N__39167),
            .I(N__39164));
    LocalMux I__8302 (
            .O(N__39164),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    CascadeMux I__8301 (
            .O(N__39161),
            .I(N__39157));
    InMux I__8300 (
            .O(N__39160),
            .I(N__39154));
    InMux I__8299 (
            .O(N__39157),
            .I(N__39151));
    LocalMux I__8298 (
            .O(N__39154),
            .I(\current_shift_inst.N_1318_i ));
    LocalMux I__8297 (
            .O(N__39151),
            .I(\current_shift_inst.N_1318_i ));
    InMux I__8296 (
            .O(N__39146),
            .I(N__39143));
    LocalMux I__8295 (
            .O(N__39143),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__8294 (
            .O(N__39140),
            .I(N__39137));
    LocalMux I__8293 (
            .O(N__39137),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__8292 (
            .O(N__39134),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__8291 (
            .O(N__39131),
            .I(N__39128));
    LocalMux I__8290 (
            .O(N__39128),
            .I(N__39124));
    InMux I__8289 (
            .O(N__39127),
            .I(N__39121));
    Span4Mux_v I__8288 (
            .O(N__39124),
            .I(N__39118));
    LocalMux I__8287 (
            .O(N__39121),
            .I(N__39115));
    Span4Mux_v I__8286 (
            .O(N__39118),
            .I(N__39110));
    Span4Mux_v I__8285 (
            .O(N__39115),
            .I(N__39107));
    InMux I__8284 (
            .O(N__39114),
            .I(N__39104));
    InMux I__8283 (
            .O(N__39113),
            .I(N__39101));
    Odrv4 I__8282 (
            .O(N__39110),
            .I(measured_delay_tr_17));
    Odrv4 I__8281 (
            .O(N__39107),
            .I(measured_delay_tr_17));
    LocalMux I__8280 (
            .O(N__39104),
            .I(measured_delay_tr_17));
    LocalMux I__8279 (
            .O(N__39101),
            .I(measured_delay_tr_17));
    CascadeMux I__8278 (
            .O(N__39092),
            .I(N__39089));
    InMux I__8277 (
            .O(N__39089),
            .I(N__39086));
    LocalMux I__8276 (
            .O(N__39086),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__8275 (
            .O(N__39083),
            .I(N__39080));
    LocalMux I__8274 (
            .O(N__39080),
            .I(N__39076));
    InMux I__8273 (
            .O(N__39079),
            .I(N__39073));
    Span4Mux_v I__8272 (
            .O(N__39076),
            .I(N__39067));
    LocalMux I__8271 (
            .O(N__39073),
            .I(N__39067));
    InMux I__8270 (
            .O(N__39072),
            .I(N__39064));
    Span4Mux_h I__8269 (
            .O(N__39067),
            .I(N__39060));
    LocalMux I__8268 (
            .O(N__39064),
            .I(N__39057));
    InMux I__8267 (
            .O(N__39063),
            .I(N__39054));
    Odrv4 I__8266 (
            .O(N__39060),
            .I(measured_delay_tr_18));
    Odrv4 I__8265 (
            .O(N__39057),
            .I(measured_delay_tr_18));
    LocalMux I__8264 (
            .O(N__39054),
            .I(measured_delay_tr_18));
    CascadeMux I__8263 (
            .O(N__39047),
            .I(N__39044));
    InMux I__8262 (
            .O(N__39044),
            .I(N__39041));
    LocalMux I__8261 (
            .O(N__39041),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CEMux I__8260 (
            .O(N__39038),
            .I(N__39033));
    CEMux I__8259 (
            .O(N__39037),
            .I(N__39030));
    CEMux I__8258 (
            .O(N__39036),
            .I(N__39027));
    LocalMux I__8257 (
            .O(N__39033),
            .I(N__39023));
    LocalMux I__8256 (
            .O(N__39030),
            .I(N__39020));
    LocalMux I__8255 (
            .O(N__39027),
            .I(N__39017));
    CEMux I__8254 (
            .O(N__39026),
            .I(N__39014));
    Odrv4 I__8253 (
            .O(N__39023),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__8252 (
            .O(N__39020),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__8251 (
            .O(N__39017),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    LocalMux I__8250 (
            .O(N__39014),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__8249 (
            .O(N__39005),
            .I(N__39002));
    InMux I__8248 (
            .O(N__39002),
            .I(N__38999));
    LocalMux I__8247 (
            .O(N__38999),
            .I(N__38996));
    Odrv4 I__8246 (
            .O(N__38996),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__8245 (
            .O(N__38993),
            .I(N__38990));
    LocalMux I__8244 (
            .O(N__38990),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__8243 (
            .O(N__38987),
            .I(N__38984));
    InMux I__8242 (
            .O(N__38984),
            .I(N__38981));
    LocalMux I__8241 (
            .O(N__38981),
            .I(N__38978));
    Odrv4 I__8240 (
            .O(N__38978),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__8239 (
            .O(N__38975),
            .I(N__38972));
    LocalMux I__8238 (
            .O(N__38972),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__8237 (
            .O(N__38969),
            .I(N__38966));
    InMux I__8236 (
            .O(N__38966),
            .I(N__38963));
    LocalMux I__8235 (
            .O(N__38963),
            .I(N__38960));
    Span4Mux_v I__8234 (
            .O(N__38960),
            .I(N__38957));
    Odrv4 I__8233 (
            .O(N__38957),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__8232 (
            .O(N__38954),
            .I(N__38951));
    LocalMux I__8231 (
            .O(N__38951),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__8230 (
            .O(N__38948),
            .I(N__38945));
    InMux I__8229 (
            .O(N__38945),
            .I(N__38942));
    LocalMux I__8228 (
            .O(N__38942),
            .I(N__38939));
    Odrv4 I__8227 (
            .O(N__38939),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__8226 (
            .O(N__38936),
            .I(N__38933));
    LocalMux I__8225 (
            .O(N__38933),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__8224 (
            .O(N__38930),
            .I(N__38927));
    InMux I__8223 (
            .O(N__38927),
            .I(N__38924));
    LocalMux I__8222 (
            .O(N__38924),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__8221 (
            .O(N__38921),
            .I(N__38918));
    LocalMux I__8220 (
            .O(N__38918),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    InMux I__8219 (
            .O(N__38915),
            .I(N__38912));
    LocalMux I__8218 (
            .O(N__38912),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__8217 (
            .O(N__38909),
            .I(N__38906));
    LocalMux I__8216 (
            .O(N__38906),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    CascadeMux I__8215 (
            .O(N__38903),
            .I(N__38900));
    InMux I__8214 (
            .O(N__38900),
            .I(N__38897));
    LocalMux I__8213 (
            .O(N__38897),
            .I(N__38894));
    Span4Mux_h I__8212 (
            .O(N__38894),
            .I(N__38891));
    Odrv4 I__8211 (
            .O(N__38891),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__8210 (
            .O(N__38888),
            .I(N__38885));
    LocalMux I__8209 (
            .O(N__38885),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    CascadeMux I__8208 (
            .O(N__38882),
            .I(N__38879));
    InMux I__8207 (
            .O(N__38879),
            .I(N__38876));
    LocalMux I__8206 (
            .O(N__38876),
            .I(N__38873));
    Odrv4 I__8205 (
            .O(N__38873),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__8204 (
            .O(N__38870),
            .I(N__38867));
    LocalMux I__8203 (
            .O(N__38867),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__8202 (
            .O(N__38864),
            .I(N__38861));
    InMux I__8201 (
            .O(N__38861),
            .I(N__38858));
    LocalMux I__8200 (
            .O(N__38858),
            .I(N__38855));
    Odrv4 I__8199 (
            .O(N__38855),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__8198 (
            .O(N__38852),
            .I(N__38849));
    LocalMux I__8197 (
            .O(N__38849),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__8196 (
            .O(N__38846),
            .I(N__38843));
    InMux I__8195 (
            .O(N__38843),
            .I(N__38840));
    LocalMux I__8194 (
            .O(N__38840),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__8193 (
            .O(N__38837),
            .I(N__38834));
    LocalMux I__8192 (
            .O(N__38834),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__8191 (
            .O(N__38831),
            .I(N__38828));
    InMux I__8190 (
            .O(N__38828),
            .I(N__38825));
    LocalMux I__8189 (
            .O(N__38825),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__8188 (
            .O(N__38822),
            .I(N__38819));
    LocalMux I__8187 (
            .O(N__38819),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__8186 (
            .O(N__38816),
            .I(N__38813));
    InMux I__8185 (
            .O(N__38813),
            .I(N__38810));
    LocalMux I__8184 (
            .O(N__38810),
            .I(N__38807));
    Odrv4 I__8183 (
            .O(N__38807),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__8182 (
            .O(N__38804),
            .I(N__38801));
    LocalMux I__8181 (
            .O(N__38801),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__8180 (
            .O(N__38798),
            .I(N__38795));
    InMux I__8179 (
            .O(N__38795),
            .I(N__38792));
    LocalMux I__8178 (
            .O(N__38792),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__8177 (
            .O(N__38789),
            .I(N__38786));
    LocalMux I__8176 (
            .O(N__38786),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__8175 (
            .O(N__38783),
            .I(N__38780));
    InMux I__8174 (
            .O(N__38780),
            .I(N__38777));
    LocalMux I__8173 (
            .O(N__38777),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__8172 (
            .O(N__38774),
            .I(N__38771));
    LocalMux I__8171 (
            .O(N__38771),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__8170 (
            .O(N__38768),
            .I(N__38765));
    InMux I__8169 (
            .O(N__38765),
            .I(N__38762));
    LocalMux I__8168 (
            .O(N__38762),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8167 (
            .O(N__38759),
            .I(N__38756));
    LocalMux I__8166 (
            .O(N__38756),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__8165 (
            .O(N__38753),
            .I(N__38750));
    LocalMux I__8164 (
            .O(N__38750),
            .I(N__38744));
    InMux I__8163 (
            .O(N__38749),
            .I(N__38741));
    CascadeMux I__8162 (
            .O(N__38748),
            .I(N__38738));
    CascadeMux I__8161 (
            .O(N__38747),
            .I(N__38735));
    Span4Mux_v I__8160 (
            .O(N__38744),
            .I(N__38730));
    LocalMux I__8159 (
            .O(N__38741),
            .I(N__38730));
    InMux I__8158 (
            .O(N__38738),
            .I(N__38727));
    InMux I__8157 (
            .O(N__38735),
            .I(N__38724));
    Odrv4 I__8156 (
            .O(N__38730),
            .I(measured_delay_tr_19));
    LocalMux I__8155 (
            .O(N__38727),
            .I(measured_delay_tr_19));
    LocalMux I__8154 (
            .O(N__38724),
            .I(measured_delay_tr_19));
    InMux I__8153 (
            .O(N__38717),
            .I(N__38714));
    LocalMux I__8152 (
            .O(N__38714),
            .I(N__38710));
    InMux I__8151 (
            .O(N__38713),
            .I(N__38707));
    Span4Mux_h I__8150 (
            .O(N__38710),
            .I(N__38701));
    LocalMux I__8149 (
            .O(N__38707),
            .I(N__38701));
    InMux I__8148 (
            .O(N__38706),
            .I(N__38698));
    Odrv4 I__8147 (
            .O(N__38701),
            .I(measured_delay_tr_12));
    LocalMux I__8146 (
            .O(N__38698),
            .I(measured_delay_tr_12));
    InMux I__8145 (
            .O(N__38693),
            .I(N__38689));
    InMux I__8144 (
            .O(N__38692),
            .I(N__38683));
    LocalMux I__8143 (
            .O(N__38689),
            .I(N__38680));
    InMux I__8142 (
            .O(N__38688),
            .I(N__38677));
    InMux I__8141 (
            .O(N__38687),
            .I(N__38672));
    InMux I__8140 (
            .O(N__38686),
            .I(N__38672));
    LocalMux I__8139 (
            .O(N__38683),
            .I(N__38669));
    Span4Mux_h I__8138 (
            .O(N__38680),
            .I(N__38664));
    LocalMux I__8137 (
            .O(N__38677),
            .I(N__38664));
    LocalMux I__8136 (
            .O(N__38672),
            .I(N__38661));
    Span4Mux_h I__8135 (
            .O(N__38669),
            .I(N__38658));
    Span4Mux_v I__8134 (
            .O(N__38664),
            .I(N__38655));
    Span4Mux_h I__8133 (
            .O(N__38661),
            .I(N__38652));
    Odrv4 I__8132 (
            .O(N__38658),
            .I(measured_delay_tr_14));
    Odrv4 I__8131 (
            .O(N__38655),
            .I(measured_delay_tr_14));
    Odrv4 I__8130 (
            .O(N__38652),
            .I(measured_delay_tr_14));
    InMux I__8129 (
            .O(N__38645),
            .I(N__38636));
    InMux I__8128 (
            .O(N__38644),
            .I(N__38636));
    InMux I__8127 (
            .O(N__38643),
            .I(N__38631));
    InMux I__8126 (
            .O(N__38642),
            .I(N__38631));
    CascadeMux I__8125 (
            .O(N__38641),
            .I(N__38628));
    LocalMux I__8124 (
            .O(N__38636),
            .I(N__38623));
    LocalMux I__8123 (
            .O(N__38631),
            .I(N__38620));
    InMux I__8122 (
            .O(N__38628),
            .I(N__38613));
    InMux I__8121 (
            .O(N__38627),
            .I(N__38613));
    InMux I__8120 (
            .O(N__38626),
            .I(N__38613));
    Span4Mux_h I__8119 (
            .O(N__38623),
            .I(N__38608));
    Span4Mux_h I__8118 (
            .O(N__38620),
            .I(N__38603));
    LocalMux I__8117 (
            .O(N__38613),
            .I(N__38603));
    InMux I__8116 (
            .O(N__38612),
            .I(N__38598));
    InMux I__8115 (
            .O(N__38611),
            .I(N__38598));
    Odrv4 I__8114 (
            .O(N__38608),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    Odrv4 I__8113 (
            .O(N__38603),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__8112 (
            .O(N__38598),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    InMux I__8111 (
            .O(N__38591),
            .I(N__38587));
    InMux I__8110 (
            .O(N__38590),
            .I(N__38584));
    LocalMux I__8109 (
            .O(N__38587),
            .I(N__38580));
    LocalMux I__8108 (
            .O(N__38584),
            .I(N__38577));
    CascadeMux I__8107 (
            .O(N__38583),
            .I(N__38574));
    Span4Mux_v I__8106 (
            .O(N__38580),
            .I(N__38571));
    Span4Mux_h I__8105 (
            .O(N__38577),
            .I(N__38568));
    InMux I__8104 (
            .O(N__38574),
            .I(N__38565));
    Odrv4 I__8103 (
            .O(N__38571),
            .I(measured_delay_tr_13));
    Odrv4 I__8102 (
            .O(N__38568),
            .I(measured_delay_tr_13));
    LocalMux I__8101 (
            .O(N__38565),
            .I(measured_delay_tr_13));
    InMux I__8100 (
            .O(N__38558),
            .I(N__38552));
    InMux I__8099 (
            .O(N__38557),
            .I(N__38552));
    LocalMux I__8098 (
            .O(N__38552),
            .I(N__38546));
    InMux I__8097 (
            .O(N__38551),
            .I(N__38542));
    InMux I__8096 (
            .O(N__38550),
            .I(N__38539));
    InMux I__8095 (
            .O(N__38549),
            .I(N__38536));
    Span4Mux_v I__8094 (
            .O(N__38546),
            .I(N__38533));
    InMux I__8093 (
            .O(N__38545),
            .I(N__38530));
    LocalMux I__8092 (
            .O(N__38542),
            .I(N__38527));
    LocalMux I__8091 (
            .O(N__38539),
            .I(N__38524));
    LocalMux I__8090 (
            .O(N__38536),
            .I(N__38521));
    Span4Mux_v I__8089 (
            .O(N__38533),
            .I(N__38516));
    LocalMux I__8088 (
            .O(N__38530),
            .I(N__38516));
    Span4Mux_v I__8087 (
            .O(N__38527),
            .I(N__38513));
    Span4Mux_h I__8086 (
            .O(N__38524),
            .I(N__38506));
    Span4Mux_v I__8085 (
            .O(N__38521),
            .I(N__38506));
    Span4Mux_h I__8084 (
            .O(N__38516),
            .I(N__38506));
    Odrv4 I__8083 (
            .O(N__38513),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    Odrv4 I__8082 (
            .O(N__38506),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    InMux I__8081 (
            .O(N__38501),
            .I(N__38492));
    InMux I__8080 (
            .O(N__38500),
            .I(N__38492));
    InMux I__8079 (
            .O(N__38499),
            .I(N__38489));
    InMux I__8078 (
            .O(N__38498),
            .I(N__38485));
    InMux I__8077 (
            .O(N__38497),
            .I(N__38482));
    LocalMux I__8076 (
            .O(N__38492),
            .I(N__38479));
    LocalMux I__8075 (
            .O(N__38489),
            .I(N__38476));
    InMux I__8074 (
            .O(N__38488),
            .I(N__38473));
    LocalMux I__8073 (
            .O(N__38485),
            .I(N__38468));
    LocalMux I__8072 (
            .O(N__38482),
            .I(N__38463));
    Span4Mux_h I__8071 (
            .O(N__38479),
            .I(N__38463));
    Span4Mux_h I__8070 (
            .O(N__38476),
            .I(N__38457));
    LocalMux I__8069 (
            .O(N__38473),
            .I(N__38457));
    InMux I__8068 (
            .O(N__38472),
            .I(N__38454));
    CascadeMux I__8067 (
            .O(N__38471),
            .I(N__38450));
    Span4Mux_v I__8066 (
            .O(N__38468),
            .I(N__38447));
    Span4Mux_v I__8065 (
            .O(N__38463),
            .I(N__38444));
    InMux I__8064 (
            .O(N__38462),
            .I(N__38441));
    Sp12to4 I__8063 (
            .O(N__38457),
            .I(N__38436));
    LocalMux I__8062 (
            .O(N__38454),
            .I(N__38436));
    InMux I__8061 (
            .O(N__38453),
            .I(N__38431));
    InMux I__8060 (
            .O(N__38450),
            .I(N__38431));
    Odrv4 I__8059 (
            .O(N__38447),
            .I(measured_delay_tr_15));
    Odrv4 I__8058 (
            .O(N__38444),
            .I(measured_delay_tr_15));
    LocalMux I__8057 (
            .O(N__38441),
            .I(measured_delay_tr_15));
    Odrv12 I__8056 (
            .O(N__38436),
            .I(measured_delay_tr_15));
    LocalMux I__8055 (
            .O(N__38431),
            .I(measured_delay_tr_15));
    CascadeMux I__8054 (
            .O(N__38420),
            .I(N__38417));
    InMux I__8053 (
            .O(N__38417),
            .I(N__38414));
    LocalMux I__8052 (
            .O(N__38414),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__8051 (
            .O(N__38411),
            .I(N__38408));
    LocalMux I__8050 (
            .O(N__38408),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__8049 (
            .O(N__38405),
            .I(N__38402));
    InMux I__8048 (
            .O(N__38402),
            .I(N__38399));
    LocalMux I__8047 (
            .O(N__38399),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__8046 (
            .O(N__38396),
            .I(N__38393));
    LocalMux I__8045 (
            .O(N__38393),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__8044 (
            .O(N__38390),
            .I(N__38387));
    InMux I__8043 (
            .O(N__38387),
            .I(N__38384));
    LocalMux I__8042 (
            .O(N__38384),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__8041 (
            .O(N__38381),
            .I(N__38378));
    LocalMux I__8040 (
            .O(N__38378),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__8039 (
            .O(N__38375),
            .I(N__38372));
    LocalMux I__8038 (
            .O(N__38372),
            .I(N__38368));
    InMux I__8037 (
            .O(N__38371),
            .I(N__38365));
    Span4Mux_h I__8036 (
            .O(N__38368),
            .I(N__38360));
    LocalMux I__8035 (
            .O(N__38365),
            .I(N__38360));
    Span4Mux_v I__8034 (
            .O(N__38360),
            .I(N__38356));
    InMux I__8033 (
            .O(N__38359),
            .I(N__38353));
    Odrv4 I__8032 (
            .O(N__38356),
            .I(measured_delay_tr_10));
    LocalMux I__8031 (
            .O(N__38353),
            .I(measured_delay_tr_10));
    CascadeMux I__8030 (
            .O(N__38348),
            .I(N__38345));
    InMux I__8029 (
            .O(N__38345),
            .I(N__38342));
    LocalMux I__8028 (
            .O(N__38342),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__8027 (
            .O(N__38339),
            .I(N__38336));
    InMux I__8026 (
            .O(N__38336),
            .I(N__38333));
    LocalMux I__8025 (
            .O(N__38333),
            .I(N__38330));
    Odrv4 I__8024 (
            .O(N__38330),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__8023 (
            .O(N__38327),
            .I(N__38324));
    InMux I__8022 (
            .O(N__38324),
            .I(N__38321));
    LocalMux I__8021 (
            .O(N__38321),
            .I(N__38318));
    Odrv4 I__8020 (
            .O(N__38318),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__8019 (
            .O(N__38315),
            .I(N__38308));
    InMux I__8018 (
            .O(N__38314),
            .I(N__38298));
    InMux I__8017 (
            .O(N__38313),
            .I(N__38298));
    InMux I__8016 (
            .O(N__38312),
            .I(N__38298));
    InMux I__8015 (
            .O(N__38311),
            .I(N__38298));
    InMux I__8014 (
            .O(N__38308),
            .I(N__38292));
    InMux I__8013 (
            .O(N__38307),
            .I(N__38292));
    LocalMux I__8012 (
            .O(N__38298),
            .I(N__38289));
    InMux I__8011 (
            .O(N__38297),
            .I(N__38286));
    LocalMux I__8010 (
            .O(N__38292),
            .I(N__38282));
    Span4Mux_h I__8009 (
            .O(N__38289),
            .I(N__38277));
    LocalMux I__8008 (
            .O(N__38286),
            .I(N__38277));
    InMux I__8007 (
            .O(N__38285),
            .I(N__38271));
    Span4Mux_v I__8006 (
            .O(N__38282),
            .I(N__38268));
    Span4Mux_v I__8005 (
            .O(N__38277),
            .I(N__38265));
    InMux I__8004 (
            .O(N__38276),
            .I(N__38258));
    InMux I__8003 (
            .O(N__38275),
            .I(N__38258));
    InMux I__8002 (
            .O(N__38274),
            .I(N__38258));
    LocalMux I__8001 (
            .O(N__38271),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    Odrv4 I__8000 (
            .O(N__38268),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    Odrv4 I__7999 (
            .O(N__38265),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__7998 (
            .O(N__38258),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    InMux I__7997 (
            .O(N__38249),
            .I(N__38245));
    InMux I__7996 (
            .O(N__38248),
            .I(N__38242));
    LocalMux I__7995 (
            .O(N__38245),
            .I(N__38236));
    LocalMux I__7994 (
            .O(N__38242),
            .I(N__38236));
    InMux I__7993 (
            .O(N__38241),
            .I(N__38233));
    Span4Mux_v I__7992 (
            .O(N__38236),
            .I(N__38230));
    LocalMux I__7991 (
            .O(N__38233),
            .I(N__38227));
    Odrv4 I__7990 (
            .O(N__38230),
            .I(measured_delay_tr_4));
    Odrv4 I__7989 (
            .O(N__38227),
            .I(measured_delay_tr_4));
    CascadeMux I__7988 (
            .O(N__38222),
            .I(N__38219));
    InMux I__7987 (
            .O(N__38219),
            .I(N__38216));
    LocalMux I__7986 (
            .O(N__38216),
            .I(N__38213));
    Odrv4 I__7985 (
            .O(N__38213),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__7984 (
            .O(N__38210),
            .I(N__38205));
    InMux I__7983 (
            .O(N__38209),
            .I(N__38202));
    InMux I__7982 (
            .O(N__38208),
            .I(N__38199));
    LocalMux I__7981 (
            .O(N__38205),
            .I(N__38196));
    LocalMux I__7980 (
            .O(N__38202),
            .I(N__38193));
    LocalMux I__7979 (
            .O(N__38199),
            .I(N__38186));
    Span4Mux_v I__7978 (
            .O(N__38196),
            .I(N__38186));
    Span4Mux_v I__7977 (
            .O(N__38193),
            .I(N__38186));
    Odrv4 I__7976 (
            .O(N__38186),
            .I(\phase_controller_inst2.stoper_tr.time_passed11 ));
    InMux I__7975 (
            .O(N__38183),
            .I(N__38178));
    InMux I__7974 (
            .O(N__38182),
            .I(N__38173));
    InMux I__7973 (
            .O(N__38181),
            .I(N__38169));
    LocalMux I__7972 (
            .O(N__38178),
            .I(N__38166));
    InMux I__7971 (
            .O(N__38177),
            .I(N__38161));
    InMux I__7970 (
            .O(N__38176),
            .I(N__38161));
    LocalMux I__7969 (
            .O(N__38173),
            .I(N__38158));
    InMux I__7968 (
            .O(N__38172),
            .I(N__38155));
    LocalMux I__7967 (
            .O(N__38169),
            .I(N__38152));
    Odrv4 I__7966 (
            .O(N__38166),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__7965 (
            .O(N__38161),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__7964 (
            .O(N__38158),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__7963 (
            .O(N__38155),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__7962 (
            .O(N__38152),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__7961 (
            .O(N__38141),
            .I(N__38138));
    LocalMux I__7960 (
            .O(N__38138),
            .I(N__38135));
    Span4Mux_s3_v I__7959 (
            .O(N__38135),
            .I(N__38132));
    Odrv4 I__7958 (
            .O(N__38132),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ));
    InMux I__7957 (
            .O(N__38129),
            .I(N__38126));
    LocalMux I__7956 (
            .O(N__38126),
            .I(N__38123));
    Span4Mux_h I__7955 (
            .O(N__38123),
            .I(N__38120));
    Odrv4 I__7954 (
            .O(N__38120),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ));
    InMux I__7953 (
            .O(N__38117),
            .I(N__38114));
    LocalMux I__7952 (
            .O(N__38114),
            .I(N__38111));
    Span4Mux_v I__7951 (
            .O(N__38111),
            .I(N__38108));
    Odrv4 I__7950 (
            .O(N__38108),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ));
    CascadeMux I__7949 (
            .O(N__38105),
            .I(N__38102));
    InMux I__7948 (
            .O(N__38102),
            .I(N__38088));
    InMux I__7947 (
            .O(N__38101),
            .I(N__38081));
    InMux I__7946 (
            .O(N__38100),
            .I(N__38081));
    InMux I__7945 (
            .O(N__38099),
            .I(N__38081));
    InMux I__7944 (
            .O(N__38098),
            .I(N__38078));
    InMux I__7943 (
            .O(N__38097),
            .I(N__38069));
    InMux I__7942 (
            .O(N__38096),
            .I(N__38069));
    InMux I__7941 (
            .O(N__38095),
            .I(N__38069));
    InMux I__7940 (
            .O(N__38094),
            .I(N__38069));
    InMux I__7939 (
            .O(N__38093),
            .I(N__38060));
    InMux I__7938 (
            .O(N__38092),
            .I(N__38060));
    InMux I__7937 (
            .O(N__38091),
            .I(N__38060));
    LocalMux I__7936 (
            .O(N__38088),
            .I(N__38053));
    LocalMux I__7935 (
            .O(N__38081),
            .I(N__38053));
    LocalMux I__7934 (
            .O(N__38078),
            .I(N__38053));
    LocalMux I__7933 (
            .O(N__38069),
            .I(N__38050));
    InMux I__7932 (
            .O(N__38068),
            .I(N__38047));
    InMux I__7931 (
            .O(N__38067),
            .I(N__38042));
    LocalMux I__7930 (
            .O(N__38060),
            .I(N__38039));
    Sp12to4 I__7929 (
            .O(N__38053),
            .I(N__38032));
    Sp12to4 I__7928 (
            .O(N__38050),
            .I(N__38032));
    LocalMux I__7927 (
            .O(N__38047),
            .I(N__38032));
    InMux I__7926 (
            .O(N__38046),
            .I(N__38027));
    InMux I__7925 (
            .O(N__38045),
            .I(N__38027));
    LocalMux I__7924 (
            .O(N__38042),
            .I(N__38022));
    Span4Mux_h I__7923 (
            .O(N__38039),
            .I(N__38022));
    Span12Mux_v I__7922 (
            .O(N__38032),
            .I(N__38019));
    LocalMux I__7921 (
            .O(N__38027),
            .I(N__38014));
    Span4Mux_v I__7920 (
            .O(N__38022),
            .I(N__38014));
    Odrv12 I__7919 (
            .O(N__38019),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    Odrv4 I__7918 (
            .O(N__38014),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    CascadeMux I__7917 (
            .O(N__38009),
            .I(N__38006));
    InMux I__7916 (
            .O(N__38006),
            .I(N__38003));
    LocalMux I__7915 (
            .O(N__38003),
            .I(\phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__7914 (
            .O(N__38000),
            .I(N__37997));
    LocalMux I__7913 (
            .O(N__37997),
            .I(N__37993));
    InMux I__7912 (
            .O(N__37996),
            .I(N__37990));
    Sp12to4 I__7911 (
            .O(N__37993),
            .I(N__37984));
    LocalMux I__7910 (
            .O(N__37990),
            .I(N__37984));
    InMux I__7909 (
            .O(N__37989),
            .I(N__37981));
    Span12Mux_v I__7908 (
            .O(N__37984),
            .I(N__37978));
    LocalMux I__7907 (
            .O(N__37981),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv12 I__7906 (
            .O(N__37978),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__7905 (
            .O(N__37973),
            .I(N__37970));
    InMux I__7904 (
            .O(N__37970),
            .I(N__37967));
    LocalMux I__7903 (
            .O(N__37967),
            .I(N__37964));
    Odrv12 I__7902 (
            .O(N__37964),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__7901 (
            .O(N__37961),
            .I(N__37958));
    LocalMux I__7900 (
            .O(N__37958),
            .I(N__37954));
    InMux I__7899 (
            .O(N__37957),
            .I(N__37951));
    Odrv4 I__7898 (
            .O(N__37954),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__7897 (
            .O(N__37951),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7896 (
            .O(N__37946),
            .I(N__37943));
    LocalMux I__7895 (
            .O(N__37943),
            .I(N__37940));
    Odrv4 I__7894 (
            .O(N__37940),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ));
    CascadeMux I__7893 (
            .O(N__37937),
            .I(N__37934));
    InMux I__7892 (
            .O(N__37934),
            .I(N__37931));
    LocalMux I__7891 (
            .O(N__37931),
            .I(N__37927));
    InMux I__7890 (
            .O(N__37930),
            .I(N__37924));
    Odrv4 I__7889 (
            .O(N__37927),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__7888 (
            .O(N__37924),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__7887 (
            .O(N__37919),
            .I(N__37916));
    LocalMux I__7886 (
            .O(N__37916),
            .I(N__37913));
    Odrv4 I__7885 (
            .O(N__37913),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__7884 (
            .O(N__37910),
            .I(N__37907));
    LocalMux I__7883 (
            .O(N__37907),
            .I(N__37903));
    InMux I__7882 (
            .O(N__37906),
            .I(N__37900));
    Odrv12 I__7881 (
            .O(N__37903),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__7880 (
            .O(N__37900),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__7879 (
            .O(N__37895),
            .I(N__37892));
    InMux I__7878 (
            .O(N__37892),
            .I(N__37889));
    LocalMux I__7877 (
            .O(N__37889),
            .I(N__37886));
    Odrv4 I__7876 (
            .O(N__37886),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__7875 (
            .O(N__37883),
            .I(N__37880));
    LocalMux I__7874 (
            .O(N__37880),
            .I(N__37877));
    Span4Mux_s1_v I__7873 (
            .O(N__37877),
            .I(N__37873));
    InMux I__7872 (
            .O(N__37876),
            .I(N__37870));
    Odrv4 I__7871 (
            .O(N__37873),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__7870 (
            .O(N__37870),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7869 (
            .O(N__37865),
            .I(N__37862));
    LocalMux I__7868 (
            .O(N__37862),
            .I(N__37859));
    Odrv12 I__7867 (
            .O(N__37859),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__7866 (
            .O(N__37856),
            .I(N__37853));
    LocalMux I__7865 (
            .O(N__37853),
            .I(N__37849));
    InMux I__7864 (
            .O(N__37852),
            .I(N__37846));
    Odrv4 I__7863 (
            .O(N__37849),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__7862 (
            .O(N__37846),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__7861 (
            .O(N__37841),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__7860 (
            .O(N__37838),
            .I(N__37835));
    InMux I__7859 (
            .O(N__37835),
            .I(N__37831));
    InMux I__7858 (
            .O(N__37834),
            .I(N__37827));
    LocalMux I__7857 (
            .O(N__37831),
            .I(N__37824));
    InMux I__7856 (
            .O(N__37830),
            .I(N__37821));
    LocalMux I__7855 (
            .O(N__37827),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__7854 (
            .O(N__37824),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__7853 (
            .O(N__37821),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__7852 (
            .O(N__37814),
            .I(N__37806));
    CascadeMux I__7851 (
            .O(N__37813),
            .I(N__37797));
    CascadeMux I__7850 (
            .O(N__37812),
            .I(N__37794));
    InMux I__7849 (
            .O(N__37811),
            .I(N__37776));
    InMux I__7848 (
            .O(N__37810),
            .I(N__37776));
    InMux I__7847 (
            .O(N__37809),
            .I(N__37776));
    LocalMux I__7846 (
            .O(N__37806),
            .I(N__37773));
    InMux I__7845 (
            .O(N__37805),
            .I(N__37760));
    InMux I__7844 (
            .O(N__37804),
            .I(N__37760));
    InMux I__7843 (
            .O(N__37803),
            .I(N__37760));
    InMux I__7842 (
            .O(N__37802),
            .I(N__37760));
    InMux I__7841 (
            .O(N__37801),
            .I(N__37760));
    InMux I__7840 (
            .O(N__37800),
            .I(N__37760));
    InMux I__7839 (
            .O(N__37797),
            .I(N__37755));
    InMux I__7838 (
            .O(N__37794),
            .I(N__37755));
    InMux I__7837 (
            .O(N__37793),
            .I(N__37746));
    InMux I__7836 (
            .O(N__37792),
            .I(N__37746));
    InMux I__7835 (
            .O(N__37791),
            .I(N__37746));
    InMux I__7834 (
            .O(N__37790),
            .I(N__37746));
    InMux I__7833 (
            .O(N__37789),
            .I(N__37739));
    InMux I__7832 (
            .O(N__37788),
            .I(N__37739));
    InMux I__7831 (
            .O(N__37787),
            .I(N__37739));
    InMux I__7830 (
            .O(N__37786),
            .I(N__37734));
    InMux I__7829 (
            .O(N__37785),
            .I(N__37734));
    CascadeMux I__7828 (
            .O(N__37784),
            .I(N__37731));
    InMux I__7827 (
            .O(N__37783),
            .I(N__37727));
    LocalMux I__7826 (
            .O(N__37776),
            .I(N__37722));
    Span4Mux_v I__7825 (
            .O(N__37773),
            .I(N__37722));
    LocalMux I__7824 (
            .O(N__37760),
            .I(N__37719));
    LocalMux I__7823 (
            .O(N__37755),
            .I(N__37710));
    LocalMux I__7822 (
            .O(N__37746),
            .I(N__37710));
    LocalMux I__7821 (
            .O(N__37739),
            .I(N__37710));
    LocalMux I__7820 (
            .O(N__37734),
            .I(N__37710));
    InMux I__7819 (
            .O(N__37731),
            .I(N__37705));
    InMux I__7818 (
            .O(N__37730),
            .I(N__37705));
    LocalMux I__7817 (
            .O(N__37727),
            .I(N__37702));
    Span4Mux_v I__7816 (
            .O(N__37722),
            .I(N__37699));
    Span4Mux_h I__7815 (
            .O(N__37719),
            .I(N__37694));
    Span4Mux_v I__7814 (
            .O(N__37710),
            .I(N__37694));
    LocalMux I__7813 (
            .O(N__37705),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__7812 (
            .O(N__37702),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__7811 (
            .O(N__37699),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__7810 (
            .O(N__37694),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__7809 (
            .O(N__37685),
            .I(N__37678));
    CascadeMux I__7808 (
            .O(N__37684),
            .I(N__37668));
    InMux I__7807 (
            .O(N__37683),
            .I(N__37656));
    InMux I__7806 (
            .O(N__37682),
            .I(N__37656));
    InMux I__7805 (
            .O(N__37681),
            .I(N__37656));
    InMux I__7804 (
            .O(N__37678),
            .I(N__37656));
    InMux I__7803 (
            .O(N__37677),
            .I(N__37653));
    CascadeMux I__7802 (
            .O(N__37676),
            .I(N__37647));
    CascadeMux I__7801 (
            .O(N__37675),
            .I(N__37644));
    CascadeMux I__7800 (
            .O(N__37674),
            .I(N__37641));
    CascadeMux I__7799 (
            .O(N__37673),
            .I(N__37638));
    CascadeMux I__7798 (
            .O(N__37672),
            .I(N__37635));
    CascadeMux I__7797 (
            .O(N__37671),
            .I(N__37632));
    InMux I__7796 (
            .O(N__37668),
            .I(N__37623));
    InMux I__7795 (
            .O(N__37667),
            .I(N__37623));
    InMux I__7794 (
            .O(N__37666),
            .I(N__37623));
    CascadeMux I__7793 (
            .O(N__37665),
            .I(N__37619));
    LocalMux I__7792 (
            .O(N__37656),
            .I(N__37613));
    LocalMux I__7791 (
            .O(N__37653),
            .I(N__37613));
    InMux I__7790 (
            .O(N__37652),
            .I(N__37600));
    InMux I__7789 (
            .O(N__37651),
            .I(N__37600));
    InMux I__7788 (
            .O(N__37650),
            .I(N__37600));
    InMux I__7787 (
            .O(N__37647),
            .I(N__37600));
    InMux I__7786 (
            .O(N__37644),
            .I(N__37600));
    InMux I__7785 (
            .O(N__37641),
            .I(N__37600));
    InMux I__7784 (
            .O(N__37638),
            .I(N__37589));
    InMux I__7783 (
            .O(N__37635),
            .I(N__37589));
    InMux I__7782 (
            .O(N__37632),
            .I(N__37589));
    InMux I__7781 (
            .O(N__37631),
            .I(N__37589));
    InMux I__7780 (
            .O(N__37630),
            .I(N__37589));
    LocalMux I__7779 (
            .O(N__37623),
            .I(N__37586));
    InMux I__7778 (
            .O(N__37622),
            .I(N__37583));
    InMux I__7777 (
            .O(N__37619),
            .I(N__37577));
    InMux I__7776 (
            .O(N__37618),
            .I(N__37577));
    Span4Mux_s2_v I__7775 (
            .O(N__37613),
            .I(N__37573));
    LocalMux I__7774 (
            .O(N__37600),
            .I(N__37570));
    LocalMux I__7773 (
            .O(N__37589),
            .I(N__37563));
    Span4Mux_v I__7772 (
            .O(N__37586),
            .I(N__37563));
    LocalMux I__7771 (
            .O(N__37583),
            .I(N__37563));
    InMux I__7770 (
            .O(N__37582),
            .I(N__37560));
    LocalMux I__7769 (
            .O(N__37577),
            .I(N__37557));
    InMux I__7768 (
            .O(N__37576),
            .I(N__37554));
    Span4Mux_h I__7767 (
            .O(N__37573),
            .I(N__37551));
    Span4Mux_h I__7766 (
            .O(N__37570),
            .I(N__37548));
    Span4Mux_h I__7765 (
            .O(N__37563),
            .I(N__37545));
    LocalMux I__7764 (
            .O(N__37560),
            .I(N__37538));
    Span4Mux_v I__7763 (
            .O(N__37557),
            .I(N__37538));
    LocalMux I__7762 (
            .O(N__37554),
            .I(N__37538));
    Odrv4 I__7761 (
            .O(N__37551),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7760 (
            .O(N__37548),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7759 (
            .O(N__37545),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7758 (
            .O(N__37538),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CascadeMux I__7757 (
            .O(N__37529),
            .I(N__37519));
    InMux I__7756 (
            .O(N__37528),
            .I(N__37500));
    InMux I__7755 (
            .O(N__37527),
            .I(N__37500));
    InMux I__7754 (
            .O(N__37526),
            .I(N__37500));
    InMux I__7753 (
            .O(N__37525),
            .I(N__37500));
    InMux I__7752 (
            .O(N__37524),
            .I(N__37500));
    InMux I__7751 (
            .O(N__37523),
            .I(N__37497));
    CascadeMux I__7750 (
            .O(N__37522),
            .I(N__37494));
    InMux I__7749 (
            .O(N__37519),
            .I(N__37483));
    InMux I__7748 (
            .O(N__37518),
            .I(N__37483));
    InMux I__7747 (
            .O(N__37517),
            .I(N__37470));
    InMux I__7746 (
            .O(N__37516),
            .I(N__37470));
    InMux I__7745 (
            .O(N__37515),
            .I(N__37470));
    InMux I__7744 (
            .O(N__37514),
            .I(N__37470));
    InMux I__7743 (
            .O(N__37513),
            .I(N__37470));
    InMux I__7742 (
            .O(N__37512),
            .I(N__37470));
    InMux I__7741 (
            .O(N__37511),
            .I(N__37467));
    LocalMux I__7740 (
            .O(N__37500),
            .I(N__37462));
    LocalMux I__7739 (
            .O(N__37497),
            .I(N__37462));
    InMux I__7738 (
            .O(N__37494),
            .I(N__37457));
    InMux I__7737 (
            .O(N__37493),
            .I(N__37457));
    InMux I__7736 (
            .O(N__37492),
            .I(N__37454));
    InMux I__7735 (
            .O(N__37491),
            .I(N__37445));
    InMux I__7734 (
            .O(N__37490),
            .I(N__37445));
    InMux I__7733 (
            .O(N__37489),
            .I(N__37445));
    InMux I__7732 (
            .O(N__37488),
            .I(N__37445));
    LocalMux I__7731 (
            .O(N__37483),
            .I(N__37442));
    LocalMux I__7730 (
            .O(N__37470),
            .I(N__37437));
    LocalMux I__7729 (
            .O(N__37467),
            .I(N__37432));
    Span4Mux_h I__7728 (
            .O(N__37462),
            .I(N__37432));
    LocalMux I__7727 (
            .O(N__37457),
            .I(N__37427));
    LocalMux I__7726 (
            .O(N__37454),
            .I(N__37427));
    LocalMux I__7725 (
            .O(N__37445),
            .I(N__37424));
    Span4Mux_s1_v I__7724 (
            .O(N__37442),
            .I(N__37421));
    InMux I__7723 (
            .O(N__37441),
            .I(N__37416));
    InMux I__7722 (
            .O(N__37440),
            .I(N__37416));
    Span4Mux_h I__7721 (
            .O(N__37437),
            .I(N__37413));
    Span4Mux_v I__7720 (
            .O(N__37432),
            .I(N__37410));
    Span4Mux_h I__7719 (
            .O(N__37427),
            .I(N__37403));
    Span4Mux_v I__7718 (
            .O(N__37424),
            .I(N__37403));
    Span4Mux_v I__7717 (
            .O(N__37421),
            .I(N__37403));
    LocalMux I__7716 (
            .O(N__37416),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__7715 (
            .O(N__37413),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__7714 (
            .O(N__37410),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__7713 (
            .O(N__37403),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__7712 (
            .O(N__37394),
            .I(N__37391));
    LocalMux I__7711 (
            .O(N__37391),
            .I(N__37388));
    Odrv4 I__7710 (
            .O(N__37388),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__7709 (
            .O(N__37385),
            .I(N__37382));
    LocalMux I__7708 (
            .O(N__37382),
            .I(N__37378));
    InMux I__7707 (
            .O(N__37381),
            .I(N__37375));
    Odrv4 I__7706 (
            .O(N__37378),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__7705 (
            .O(N__37375),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7704 (
            .O(N__37370),
            .I(N__37366));
    InMux I__7703 (
            .O(N__37369),
            .I(N__37363));
    LocalMux I__7702 (
            .O(N__37366),
            .I(N__37360));
    LocalMux I__7701 (
            .O(N__37363),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv12 I__7700 (
            .O(N__37360),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__7699 (
            .O(N__37355),
            .I(N__37352));
    InMux I__7698 (
            .O(N__37352),
            .I(N__37349));
    LocalMux I__7697 (
            .O(N__37349),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__7696 (
            .O(N__37346),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__7695 (
            .O(N__37343),
            .I(N__37340));
    LocalMux I__7694 (
            .O(N__37340),
            .I(N__37336));
    InMux I__7693 (
            .O(N__37339),
            .I(N__37333));
    Span4Mux_v I__7692 (
            .O(N__37336),
            .I(N__37330));
    LocalMux I__7691 (
            .O(N__37333),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__7690 (
            .O(N__37330),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__7689 (
            .O(N__37325),
            .I(N__37322));
    LocalMux I__7688 (
            .O(N__37322),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__7687 (
            .O(N__37319),
            .I(bfn_15_4_0_));
    InMux I__7686 (
            .O(N__37316),
            .I(N__37312));
    InMux I__7685 (
            .O(N__37315),
            .I(N__37309));
    LocalMux I__7684 (
            .O(N__37312),
            .I(N__37306));
    LocalMux I__7683 (
            .O(N__37309),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv12 I__7682 (
            .O(N__37306),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__7681 (
            .O(N__37301),
            .I(N__37298));
    LocalMux I__7680 (
            .O(N__37298),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__7679 (
            .O(N__37295),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__7678 (
            .O(N__37292),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__7677 (
            .O(N__37289),
            .I(N__37286));
    LocalMux I__7676 (
            .O(N__37286),
            .I(N__37283));
    Span4Mux_h I__7675 (
            .O(N__37283),
            .I(N__37280));
    Odrv4 I__7674 (
            .O(N__37280),
            .I(\delay_measurement_inst.delay_tr_timer.N_290 ));
    InMux I__7673 (
            .O(N__37277),
            .I(N__37266));
    InMux I__7672 (
            .O(N__37276),
            .I(N__37266));
    InMux I__7671 (
            .O(N__37275),
            .I(N__37266));
    InMux I__7670 (
            .O(N__37274),
            .I(N__37263));
    InMux I__7669 (
            .O(N__37273),
            .I(N__37258));
    LocalMux I__7668 (
            .O(N__37266),
            .I(N__37254));
    LocalMux I__7667 (
            .O(N__37263),
            .I(N__37251));
    InMux I__7666 (
            .O(N__37262),
            .I(N__37246));
    InMux I__7665 (
            .O(N__37261),
            .I(N__37246));
    LocalMux I__7664 (
            .O(N__37258),
            .I(N__37242));
    InMux I__7663 (
            .O(N__37257),
            .I(N__37239));
    Span4Mux_v I__7662 (
            .O(N__37254),
            .I(N__37232));
    Span4Mux_v I__7661 (
            .O(N__37251),
            .I(N__37232));
    LocalMux I__7660 (
            .O(N__37246),
            .I(N__37232));
    InMux I__7659 (
            .O(N__37245),
            .I(N__37229));
    Odrv4 I__7658 (
            .O(N__37242),
            .I(\delay_measurement_inst.N_325 ));
    LocalMux I__7657 (
            .O(N__37239),
            .I(\delay_measurement_inst.N_325 ));
    Odrv4 I__7656 (
            .O(N__37232),
            .I(\delay_measurement_inst.N_325 ));
    LocalMux I__7655 (
            .O(N__37229),
            .I(\delay_measurement_inst.N_325 ));
    InMux I__7654 (
            .O(N__37220),
            .I(N__37217));
    LocalMux I__7653 (
            .O(N__37217),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__7652 (
            .O(N__37214),
            .I(N__37211));
    LocalMux I__7651 (
            .O(N__37211),
            .I(N__37207));
    InMux I__7650 (
            .O(N__37210),
            .I(N__37204));
    Span4Mux_v I__7649 (
            .O(N__37207),
            .I(N__37201));
    LocalMux I__7648 (
            .O(N__37204),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__7647 (
            .O(N__37201),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__7646 (
            .O(N__37196),
            .I(N__37193));
    InMux I__7645 (
            .O(N__37193),
            .I(N__37190));
    LocalMux I__7644 (
            .O(N__37190),
            .I(N__37187));
    Odrv4 I__7643 (
            .O(N__37187),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__7642 (
            .O(N__37184),
            .I(N__37181));
    LocalMux I__7641 (
            .O(N__37181),
            .I(N__37177));
    InMux I__7640 (
            .O(N__37180),
            .I(N__37174));
    Odrv4 I__7639 (
            .O(N__37177),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__7638 (
            .O(N__37174),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__7637 (
            .O(N__37169),
            .I(N__37166));
    LocalMux I__7636 (
            .O(N__37166),
            .I(N__37162));
    InMux I__7635 (
            .O(N__37165),
            .I(N__37159));
    Span4Mux_v I__7634 (
            .O(N__37162),
            .I(N__37156));
    LocalMux I__7633 (
            .O(N__37159),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__7632 (
            .O(N__37156),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__7631 (
            .O(N__37151),
            .I(N__37148));
    LocalMux I__7630 (
            .O(N__37148),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__7629 (
            .O(N__37145),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__7628 (
            .O(N__37142),
            .I(N__37138));
    InMux I__7627 (
            .O(N__37141),
            .I(N__37135));
    LocalMux I__7626 (
            .O(N__37138),
            .I(N__37132));
    LocalMux I__7625 (
            .O(N__37135),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__7624 (
            .O(N__37132),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__7623 (
            .O(N__37127),
            .I(N__37124));
    LocalMux I__7622 (
            .O(N__37124),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__7621 (
            .O(N__37121),
            .I(bfn_15_3_0_));
    InMux I__7620 (
            .O(N__37118),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__7619 (
            .O(N__37115),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__7618 (
            .O(N__37112),
            .I(N__37108));
    InMux I__7617 (
            .O(N__37111),
            .I(N__37105));
    LocalMux I__7616 (
            .O(N__37108),
            .I(N__37102));
    LocalMux I__7615 (
            .O(N__37105),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv12 I__7614 (
            .O(N__37102),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__7613 (
            .O(N__37097),
            .I(N__37094));
    InMux I__7612 (
            .O(N__37094),
            .I(N__37091));
    LocalMux I__7611 (
            .O(N__37091),
            .I(N__37088));
    Odrv12 I__7610 (
            .O(N__37088),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__7609 (
            .O(N__37085),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__7608 (
            .O(N__37082),
            .I(N__37078));
    InMux I__7607 (
            .O(N__37081),
            .I(N__37075));
    LocalMux I__7606 (
            .O(N__37078),
            .I(N__37072));
    LocalMux I__7605 (
            .O(N__37075),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv12 I__7604 (
            .O(N__37072),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__7603 (
            .O(N__37067),
            .I(N__37064));
    LocalMux I__7602 (
            .O(N__37064),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__7601 (
            .O(N__37061),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__7600 (
            .O(N__37058),
            .I(N__37054));
    InMux I__7599 (
            .O(N__37057),
            .I(N__37051));
    LocalMux I__7598 (
            .O(N__37054),
            .I(N__37048));
    LocalMux I__7597 (
            .O(N__37051),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__7596 (
            .O(N__37048),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__7595 (
            .O(N__37043),
            .I(N__37040));
    LocalMux I__7594 (
            .O(N__37040),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__7593 (
            .O(N__37037),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__7592 (
            .O(N__37034),
            .I(N__37031));
    LocalMux I__7591 (
            .O(N__37031),
            .I(N__37027));
    InMux I__7590 (
            .O(N__37030),
            .I(N__37024));
    Span4Mux_v I__7589 (
            .O(N__37027),
            .I(N__37021));
    LocalMux I__7588 (
            .O(N__37024),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__7587 (
            .O(N__37021),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__7586 (
            .O(N__37016),
            .I(N__37013));
    InMux I__7585 (
            .O(N__37013),
            .I(N__37010));
    LocalMux I__7584 (
            .O(N__37010),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__7583 (
            .O(N__37007),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__7582 (
            .O(N__37004),
            .I(N__36998));
    InMux I__7581 (
            .O(N__37003),
            .I(N__36993));
    InMux I__7580 (
            .O(N__37002),
            .I(N__36993));
    InMux I__7579 (
            .O(N__37001),
            .I(N__36990));
    LocalMux I__7578 (
            .O(N__36998),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7577 (
            .O(N__36993),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7576 (
            .O(N__36990),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__7575 (
            .O(N__36983),
            .I(N__36975));
    InMux I__7574 (
            .O(N__36982),
            .I(N__36975));
    InMux I__7573 (
            .O(N__36981),
            .I(N__36972));
    InMux I__7572 (
            .O(N__36980),
            .I(N__36969));
    LocalMux I__7571 (
            .O(N__36975),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7570 (
            .O(N__36972),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7569 (
            .O(N__36969),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__7568 (
            .O(N__36962),
            .I(N__36959));
    LocalMux I__7567 (
            .O(N__36959),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__7566 (
            .O(N__36956),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__7565 (
            .O(N__36953),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__7564 (
            .O(N__36950),
            .I(N__36946));
    InMux I__7563 (
            .O(N__36949),
            .I(N__36943));
    LocalMux I__7562 (
            .O(N__36946),
            .I(N__36940));
    LocalMux I__7561 (
            .O(N__36943),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__7560 (
            .O(N__36940),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__7559 (
            .O(N__36935),
            .I(N__36932));
    LocalMux I__7558 (
            .O(N__36932),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__7557 (
            .O(N__36929),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__7556 (
            .O(N__36926),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__7555 (
            .O(N__36923),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__7554 (
            .O(N__36920),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__7553 (
            .O(N__36917),
            .I(N__36913));
    InMux I__7552 (
            .O(N__36916),
            .I(N__36910));
    LocalMux I__7551 (
            .O(N__36913),
            .I(N__36907));
    LocalMux I__7550 (
            .O(N__36910),
            .I(N__36904));
    Span4Mux_v I__7549 (
            .O(N__36907),
            .I(N__36900));
    Span4Mux_h I__7548 (
            .O(N__36904),
            .I(N__36897));
    InMux I__7547 (
            .O(N__36903),
            .I(N__36894));
    Odrv4 I__7546 (
            .O(N__36900),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    Odrv4 I__7545 (
            .O(N__36897),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    LocalMux I__7544 (
            .O(N__36894),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    CascadeMux I__7543 (
            .O(N__36887),
            .I(N__36884));
    InMux I__7542 (
            .O(N__36884),
            .I(N__36881));
    LocalMux I__7541 (
            .O(N__36881),
            .I(N__36878));
    Span4Mux_v I__7540 (
            .O(N__36878),
            .I(N__36875));
    Odrv4 I__7539 (
            .O(N__36875),
            .I(\phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa ));
    CascadeMux I__7538 (
            .O(N__36872),
            .I(N__36869));
    InMux I__7537 (
            .O(N__36869),
            .I(N__36865));
    InMux I__7536 (
            .O(N__36868),
            .I(N__36862));
    LocalMux I__7535 (
            .O(N__36865),
            .I(N__36857));
    LocalMux I__7534 (
            .O(N__36862),
            .I(N__36854));
    InMux I__7533 (
            .O(N__36861),
            .I(N__36851));
    InMux I__7532 (
            .O(N__36860),
            .I(N__36846));
    Span4Mux_v I__7531 (
            .O(N__36857),
            .I(N__36843));
    Span4Mux_v I__7530 (
            .O(N__36854),
            .I(N__36840));
    LocalMux I__7529 (
            .O(N__36851),
            .I(N__36837));
    InMux I__7528 (
            .O(N__36850),
            .I(N__36834));
    InMux I__7527 (
            .O(N__36849),
            .I(N__36831));
    LocalMux I__7526 (
            .O(N__36846),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__7525 (
            .O(N__36843),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__7524 (
            .O(N__36840),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__7523 (
            .O(N__36837),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__7522 (
            .O(N__36834),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__7521 (
            .O(N__36831),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__7520 (
            .O(N__36818),
            .I(N__36815));
    LocalMux I__7519 (
            .O(N__36815),
            .I(N__36812));
    Span4Mux_h I__7518 (
            .O(N__36812),
            .I(N__36809));
    Span4Mux_h I__7517 (
            .O(N__36809),
            .I(N__36803));
    InMux I__7516 (
            .O(N__36808),
            .I(N__36798));
    InMux I__7515 (
            .O(N__36807),
            .I(N__36798));
    InMux I__7514 (
            .O(N__36806),
            .I(N__36795));
    Sp12to4 I__7513 (
            .O(N__36803),
            .I(N__36790));
    LocalMux I__7512 (
            .O(N__36798),
            .I(N__36790));
    LocalMux I__7511 (
            .O(N__36795),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__7510 (
            .O(N__36790),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__7509 (
            .O(N__36785),
            .I(N__36782));
    LocalMux I__7508 (
            .O(N__36782),
            .I(N__36779));
    Odrv12 I__7507 (
            .O(N__36779),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__7506 (
            .O(N__36776),
            .I(N__36773));
    LocalMux I__7505 (
            .O(N__36773),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__7504 (
            .O(N__36770),
            .I(N__36767));
    LocalMux I__7503 (
            .O(N__36767),
            .I(N__36764));
    Span12Mux_v I__7502 (
            .O(N__36764),
            .I(N__36761));
    Odrv12 I__7501 (
            .O(N__36761),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__7500 (
            .O(N__36758),
            .I(N__36755));
    LocalMux I__7499 (
            .O(N__36755),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__7498 (
            .O(N__36752),
            .I(N__36749));
    LocalMux I__7497 (
            .O(N__36749),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__7496 (
            .O(N__36746),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__7495 (
            .O(N__36743),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__7494 (
            .O(N__36740),
            .I(N__36737));
    LocalMux I__7493 (
            .O(N__36737),
            .I(N__36734));
    Span12Mux_h I__7492 (
            .O(N__36734),
            .I(N__36731));
    Odrv12 I__7491 (
            .O(N__36731),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__7490 (
            .O(N__36728),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__7489 (
            .O(N__36725),
            .I(N__36722));
    LocalMux I__7488 (
            .O(N__36722),
            .I(N__36719));
    Span4Mux_h I__7487 (
            .O(N__36719),
            .I(N__36716));
    Span4Mux_v I__7486 (
            .O(N__36716),
            .I(N__36713));
    Span4Mux_h I__7485 (
            .O(N__36713),
            .I(N__36710));
    Odrv4 I__7484 (
            .O(N__36710),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__7483 (
            .O(N__36707),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__7482 (
            .O(N__36704),
            .I(N__36701));
    LocalMux I__7481 (
            .O(N__36701),
            .I(N__36698));
    Span4Mux_h I__7480 (
            .O(N__36698),
            .I(N__36695));
    Odrv4 I__7479 (
            .O(N__36695),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__7478 (
            .O(N__36692),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__7477 (
            .O(N__36689),
            .I(N__36686));
    LocalMux I__7476 (
            .O(N__36686),
            .I(N__36683));
    Span4Mux_h I__7475 (
            .O(N__36683),
            .I(N__36680));
    Span4Mux_v I__7474 (
            .O(N__36680),
            .I(N__36677));
    Span4Mux_h I__7473 (
            .O(N__36677),
            .I(N__36674));
    Odrv4 I__7472 (
            .O(N__36674),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__7471 (
            .O(N__36671),
            .I(bfn_14_17_0_));
    InMux I__7470 (
            .O(N__36668),
            .I(N__36665));
    LocalMux I__7469 (
            .O(N__36665),
            .I(N__36662));
    Odrv4 I__7468 (
            .O(N__36662),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__7467 (
            .O(N__36659),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__7466 (
            .O(N__36656),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__7465 (
            .O(N__36653),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__7464 (
            .O(N__36650),
            .I(N__36647));
    LocalMux I__7463 (
            .O(N__36647),
            .I(N__36643));
    InMux I__7462 (
            .O(N__36646),
            .I(N__36640));
    Span4Mux_v I__7461 (
            .O(N__36643),
            .I(N__36635));
    LocalMux I__7460 (
            .O(N__36640),
            .I(N__36635));
    Span4Mux_v I__7459 (
            .O(N__36635),
            .I(N__36632));
    Odrv4 I__7458 (
            .O(N__36632),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    CascadeMux I__7457 (
            .O(N__36629),
            .I(N__36623));
    CascadeMux I__7456 (
            .O(N__36628),
            .I(N__36616));
    CascadeMux I__7455 (
            .O(N__36627),
            .I(N__36613));
    CascadeMux I__7454 (
            .O(N__36626),
            .I(N__36610));
    InMux I__7453 (
            .O(N__36623),
            .I(N__36598));
    InMux I__7452 (
            .O(N__36622),
            .I(N__36583));
    InMux I__7451 (
            .O(N__36621),
            .I(N__36583));
    InMux I__7450 (
            .O(N__36620),
            .I(N__36583));
    InMux I__7449 (
            .O(N__36619),
            .I(N__36583));
    InMux I__7448 (
            .O(N__36616),
            .I(N__36583));
    InMux I__7447 (
            .O(N__36613),
            .I(N__36583));
    InMux I__7446 (
            .O(N__36610),
            .I(N__36583));
    CascadeMux I__7445 (
            .O(N__36609),
            .I(N__36580));
    InMux I__7444 (
            .O(N__36608),
            .I(N__36576));
    InMux I__7443 (
            .O(N__36607),
            .I(N__36573));
    InMux I__7442 (
            .O(N__36606),
            .I(N__36570));
    CascadeMux I__7441 (
            .O(N__36605),
            .I(N__36567));
    CascadeMux I__7440 (
            .O(N__36604),
            .I(N__36563));
    CascadeMux I__7439 (
            .O(N__36603),
            .I(N__36560));
    CascadeMux I__7438 (
            .O(N__36602),
            .I(N__36557));
    CascadeMux I__7437 (
            .O(N__36601),
            .I(N__36554));
    LocalMux I__7436 (
            .O(N__36598),
            .I(N__36544));
    LocalMux I__7435 (
            .O(N__36583),
            .I(N__36544));
    InMux I__7434 (
            .O(N__36580),
            .I(N__36539));
    InMux I__7433 (
            .O(N__36579),
            .I(N__36539));
    LocalMux I__7432 (
            .O(N__36576),
            .I(N__36536));
    LocalMux I__7431 (
            .O(N__36573),
            .I(N__36533));
    LocalMux I__7430 (
            .O(N__36570),
            .I(N__36530));
    InMux I__7429 (
            .O(N__36567),
            .I(N__36527));
    InMux I__7428 (
            .O(N__36566),
            .I(N__36510));
    InMux I__7427 (
            .O(N__36563),
            .I(N__36510));
    InMux I__7426 (
            .O(N__36560),
            .I(N__36510));
    InMux I__7425 (
            .O(N__36557),
            .I(N__36510));
    InMux I__7424 (
            .O(N__36554),
            .I(N__36510));
    InMux I__7423 (
            .O(N__36553),
            .I(N__36510));
    InMux I__7422 (
            .O(N__36552),
            .I(N__36510));
    InMux I__7421 (
            .O(N__36551),
            .I(N__36510));
    InMux I__7420 (
            .O(N__36550),
            .I(N__36505));
    InMux I__7419 (
            .O(N__36549),
            .I(N__36505));
    Span4Mux_v I__7418 (
            .O(N__36544),
            .I(N__36502));
    LocalMux I__7417 (
            .O(N__36539),
            .I(N__36493));
    Span4Mux_v I__7416 (
            .O(N__36536),
            .I(N__36493));
    Span4Mux_v I__7415 (
            .O(N__36533),
            .I(N__36493));
    Span4Mux_h I__7414 (
            .O(N__36530),
            .I(N__36493));
    LocalMux I__7413 (
            .O(N__36527),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__7412 (
            .O(N__36510),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__7411 (
            .O(N__36505),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__7410 (
            .O(N__36502),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__7409 (
            .O(N__36493),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__7408 (
            .O(N__36482),
            .I(N__36460));
    CascadeMux I__7407 (
            .O(N__36481),
            .I(N__36456));
    CascadeMux I__7406 (
            .O(N__36480),
            .I(N__36453));
    CascadeMux I__7405 (
            .O(N__36479),
            .I(N__36450));
    CascadeMux I__7404 (
            .O(N__36478),
            .I(N__36447));
    InMux I__7403 (
            .O(N__36477),
            .I(N__36443));
    InMux I__7402 (
            .O(N__36476),
            .I(N__36440));
    InMux I__7401 (
            .O(N__36475),
            .I(N__36431));
    InMux I__7400 (
            .O(N__36474),
            .I(N__36431));
    InMux I__7399 (
            .O(N__36473),
            .I(N__36431));
    InMux I__7398 (
            .O(N__36472),
            .I(N__36431));
    InMux I__7397 (
            .O(N__36471),
            .I(N__36428));
    InMux I__7396 (
            .O(N__36470),
            .I(N__36412));
    InMux I__7395 (
            .O(N__36469),
            .I(N__36412));
    InMux I__7394 (
            .O(N__36468),
            .I(N__36412));
    InMux I__7393 (
            .O(N__36467),
            .I(N__36412));
    InMux I__7392 (
            .O(N__36466),
            .I(N__36412));
    InMux I__7391 (
            .O(N__36465),
            .I(N__36412));
    InMux I__7390 (
            .O(N__36464),
            .I(N__36412));
    InMux I__7389 (
            .O(N__36463),
            .I(N__36409));
    InMux I__7388 (
            .O(N__36460),
            .I(N__36406));
    InMux I__7387 (
            .O(N__36459),
            .I(N__36403));
    InMux I__7386 (
            .O(N__36456),
            .I(N__36394));
    InMux I__7385 (
            .O(N__36453),
            .I(N__36394));
    InMux I__7384 (
            .O(N__36450),
            .I(N__36394));
    InMux I__7383 (
            .O(N__36447),
            .I(N__36394));
    InMux I__7382 (
            .O(N__36446),
            .I(N__36391));
    LocalMux I__7381 (
            .O(N__36443),
            .I(N__36388));
    LocalMux I__7380 (
            .O(N__36440),
            .I(N__36385));
    LocalMux I__7379 (
            .O(N__36431),
            .I(N__36380));
    LocalMux I__7378 (
            .O(N__36428),
            .I(N__36380));
    InMux I__7377 (
            .O(N__36427),
            .I(N__36377));
    LocalMux I__7376 (
            .O(N__36412),
            .I(N__36373));
    LocalMux I__7375 (
            .O(N__36409),
            .I(N__36366));
    LocalMux I__7374 (
            .O(N__36406),
            .I(N__36366));
    LocalMux I__7373 (
            .O(N__36403),
            .I(N__36366));
    LocalMux I__7372 (
            .O(N__36394),
            .I(N__36353));
    LocalMux I__7371 (
            .O(N__36391),
            .I(N__36353));
    Span4Mux_h I__7370 (
            .O(N__36388),
            .I(N__36353));
    Span4Mux_v I__7369 (
            .O(N__36385),
            .I(N__36353));
    Span4Mux_h I__7368 (
            .O(N__36380),
            .I(N__36353));
    LocalMux I__7367 (
            .O(N__36377),
            .I(N__36353));
    InMux I__7366 (
            .O(N__36376),
            .I(N__36350));
    Span4Mux_v I__7365 (
            .O(N__36373),
            .I(N__36347));
    Span4Mux_v I__7364 (
            .O(N__36366),
            .I(N__36344));
    Span4Mux_v I__7363 (
            .O(N__36353),
            .I(N__36341));
    LocalMux I__7362 (
            .O(N__36350),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__7361 (
            .O(N__36347),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__7360 (
            .O(N__36344),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__7359 (
            .O(N__36341),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__7358 (
            .O(N__36332),
            .I(N__36312));
    InMux I__7357 (
            .O(N__36331),
            .I(N__36297));
    InMux I__7356 (
            .O(N__36330),
            .I(N__36297));
    InMux I__7355 (
            .O(N__36329),
            .I(N__36297));
    InMux I__7354 (
            .O(N__36328),
            .I(N__36297));
    InMux I__7353 (
            .O(N__36327),
            .I(N__36297));
    InMux I__7352 (
            .O(N__36326),
            .I(N__36297));
    InMux I__7351 (
            .O(N__36325),
            .I(N__36297));
    InMux I__7350 (
            .O(N__36324),
            .I(N__36293));
    InMux I__7349 (
            .O(N__36323),
            .I(N__36290));
    InMux I__7348 (
            .O(N__36322),
            .I(N__36270));
    InMux I__7347 (
            .O(N__36321),
            .I(N__36270));
    InMux I__7346 (
            .O(N__36320),
            .I(N__36270));
    InMux I__7345 (
            .O(N__36319),
            .I(N__36270));
    InMux I__7344 (
            .O(N__36318),
            .I(N__36270));
    InMux I__7343 (
            .O(N__36317),
            .I(N__36270));
    InMux I__7342 (
            .O(N__36316),
            .I(N__36270));
    InMux I__7341 (
            .O(N__36315),
            .I(N__36270));
    LocalMux I__7340 (
            .O(N__36312),
            .I(N__36267));
    LocalMux I__7339 (
            .O(N__36297),
            .I(N__36264));
    InMux I__7338 (
            .O(N__36296),
            .I(N__36261));
    LocalMux I__7337 (
            .O(N__36293),
            .I(N__36258));
    LocalMux I__7336 (
            .O(N__36290),
            .I(N__36255));
    InMux I__7335 (
            .O(N__36289),
            .I(N__36250));
    InMux I__7334 (
            .O(N__36288),
            .I(N__36245));
    InMux I__7333 (
            .O(N__36287),
            .I(N__36245));
    LocalMux I__7332 (
            .O(N__36270),
            .I(N__36238));
    Span4Mux_v I__7331 (
            .O(N__36267),
            .I(N__36238));
    Span4Mux_h I__7330 (
            .O(N__36264),
            .I(N__36238));
    LocalMux I__7329 (
            .O(N__36261),
            .I(N__36235));
    Span4Mux_h I__7328 (
            .O(N__36258),
            .I(N__36230));
    Span4Mux_h I__7327 (
            .O(N__36255),
            .I(N__36230));
    InMux I__7326 (
            .O(N__36254),
            .I(N__36225));
    InMux I__7325 (
            .O(N__36253),
            .I(N__36225));
    LocalMux I__7324 (
            .O(N__36250),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__7323 (
            .O(N__36245),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__7322 (
            .O(N__36238),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__7321 (
            .O(N__36235),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__7320 (
            .O(N__36230),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__7319 (
            .O(N__36225),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__7318 (
            .O(N__36212),
            .I(N__36209));
    LocalMux I__7317 (
            .O(N__36209),
            .I(N__36202));
    InMux I__7316 (
            .O(N__36208),
            .I(N__36199));
    CascadeMux I__7315 (
            .O(N__36207),
            .I(N__36196));
    InMux I__7314 (
            .O(N__36206),
            .I(N__36193));
    CascadeMux I__7313 (
            .O(N__36205),
            .I(N__36190));
    Span4Mux_v I__7312 (
            .O(N__36202),
            .I(N__36187));
    LocalMux I__7311 (
            .O(N__36199),
            .I(N__36184));
    InMux I__7310 (
            .O(N__36196),
            .I(N__36181));
    LocalMux I__7309 (
            .O(N__36193),
            .I(N__36178));
    InMux I__7308 (
            .O(N__36190),
            .I(N__36175));
    Span4Mux_v I__7307 (
            .O(N__36187),
            .I(N__36172));
    Span4Mux_h I__7306 (
            .O(N__36184),
            .I(N__36169));
    LocalMux I__7305 (
            .O(N__36181),
            .I(N__36164));
    Span4Mux_h I__7304 (
            .O(N__36178),
            .I(N__36164));
    LocalMux I__7303 (
            .O(N__36175),
            .I(measured_delay_hc_31));
    Odrv4 I__7302 (
            .O(N__36172),
            .I(measured_delay_hc_31));
    Odrv4 I__7301 (
            .O(N__36169),
            .I(measured_delay_hc_31));
    Odrv4 I__7300 (
            .O(N__36164),
            .I(measured_delay_hc_31));
    InMux I__7299 (
            .O(N__36155),
            .I(N__36152));
    LocalMux I__7298 (
            .O(N__36152),
            .I(N__36149));
    Span4Mux_h I__7297 (
            .O(N__36149),
            .I(N__36144));
    InMux I__7296 (
            .O(N__36148),
            .I(N__36141));
    InMux I__7295 (
            .O(N__36147),
            .I(N__36138));
    Odrv4 I__7294 (
            .O(N__36144),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    LocalMux I__7293 (
            .O(N__36141),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    LocalMux I__7292 (
            .O(N__36138),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    InMux I__7291 (
            .O(N__36131),
            .I(N__36127));
    InMux I__7290 (
            .O(N__36130),
            .I(N__36124));
    LocalMux I__7289 (
            .O(N__36127),
            .I(N__36117));
    LocalMux I__7288 (
            .O(N__36124),
            .I(N__36117));
    InMux I__7287 (
            .O(N__36123),
            .I(N__36114));
    InMux I__7286 (
            .O(N__36122),
            .I(N__36111));
    Span4Mux_v I__7285 (
            .O(N__36117),
            .I(N__36108));
    LocalMux I__7284 (
            .O(N__36114),
            .I(N__36105));
    LocalMux I__7283 (
            .O(N__36111),
            .I(N__36102));
    Span4Mux_v I__7282 (
            .O(N__36108),
            .I(N__36099));
    Span4Mux_h I__7281 (
            .O(N__36105),
            .I(N__36096));
    Odrv12 I__7280 (
            .O(N__36102),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ));
    Odrv4 I__7279 (
            .O(N__36099),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ));
    Odrv4 I__7278 (
            .O(N__36096),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ));
    CascadeMux I__7277 (
            .O(N__36089),
            .I(N__36086));
    InMux I__7276 (
            .O(N__36086),
            .I(N__36083));
    LocalMux I__7275 (
            .O(N__36083),
            .I(N__36080));
    Odrv4 I__7274 (
            .O(N__36080),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    CEMux I__7273 (
            .O(N__36077),
            .I(N__36072));
    CEMux I__7272 (
            .O(N__36076),
            .I(N__36069));
    CEMux I__7271 (
            .O(N__36075),
            .I(N__36066));
    LocalMux I__7270 (
            .O(N__36072),
            .I(N__36063));
    LocalMux I__7269 (
            .O(N__36069),
            .I(N__36059));
    LocalMux I__7268 (
            .O(N__36066),
            .I(N__36056));
    Span4Mux_v I__7267 (
            .O(N__36063),
            .I(N__36053));
    CEMux I__7266 (
            .O(N__36062),
            .I(N__36050));
    Span4Mux_v I__7265 (
            .O(N__36059),
            .I(N__36047));
    Span4Mux_h I__7264 (
            .O(N__36056),
            .I(N__36044));
    Sp12to4 I__7263 (
            .O(N__36053),
            .I(N__36039));
    LocalMux I__7262 (
            .O(N__36050),
            .I(N__36039));
    Span4Mux_h I__7261 (
            .O(N__36047),
            .I(N__36036));
    Odrv4 I__7260 (
            .O(N__36044),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv12 I__7259 (
            .O(N__36039),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__7258 (
            .O(N__36036),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__7257 (
            .O(N__36029),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__7256 (
            .O(N__36026),
            .I(N__36023));
    LocalMux I__7255 (
            .O(N__36023),
            .I(N__36020));
    Span4Mux_h I__7254 (
            .O(N__36020),
            .I(N__36017));
    Odrv4 I__7253 (
            .O(N__36017),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ));
    InMux I__7252 (
            .O(N__36014),
            .I(N__36010));
    InMux I__7251 (
            .O(N__36013),
            .I(N__36007));
    LocalMux I__7250 (
            .O(N__36010),
            .I(N__36004));
    LocalMux I__7249 (
            .O(N__36007),
            .I(N__36001));
    Span4Mux_v I__7248 (
            .O(N__36004),
            .I(N__35998));
    Span12Mux_v I__7247 (
            .O(N__36001),
            .I(N__35995));
    Span4Mux_v I__7246 (
            .O(N__35998),
            .I(N__35992));
    Odrv12 I__7245 (
            .O(N__35995),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    Odrv4 I__7244 (
            .O(N__35992),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__7243 (
            .O(N__35987),
            .I(N__35984));
    LocalMux I__7242 (
            .O(N__35984),
            .I(N__35981));
    Span4Mux_v I__7241 (
            .O(N__35981),
            .I(N__35978));
    Odrv4 I__7240 (
            .O(N__35978),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__7239 (
            .O(N__35975),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__7238 (
            .O(N__35972),
            .I(N__35969));
    LocalMux I__7237 (
            .O(N__35969),
            .I(N__35966));
    Span4Mux_h I__7236 (
            .O(N__35966),
            .I(N__35963));
    Span4Mux_v I__7235 (
            .O(N__35963),
            .I(N__35960));
    Span4Mux_h I__7234 (
            .O(N__35960),
            .I(N__35957));
    Odrv4 I__7233 (
            .O(N__35957),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__7232 (
            .O(N__35954),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__7231 (
            .O(N__35951),
            .I(N__35948));
    LocalMux I__7230 (
            .O(N__35948),
            .I(N__35945));
    Span4Mux_v I__7229 (
            .O(N__35945),
            .I(N__35942));
    Odrv4 I__7228 (
            .O(N__35942),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__7227 (
            .O(N__35939),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__7226 (
            .O(N__35936),
            .I(N__35933));
    LocalMux I__7225 (
            .O(N__35933),
            .I(N__35930));
    Odrv4 I__7224 (
            .O(N__35930),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    CEMux I__7223 (
            .O(N__35927),
            .I(N__35924));
    LocalMux I__7222 (
            .O(N__35924),
            .I(N__35921));
    Span4Mux_v I__7221 (
            .O(N__35921),
            .I(N__35917));
    CEMux I__7220 (
            .O(N__35920),
            .I(N__35914));
    Span4Mux_v I__7219 (
            .O(N__35917),
            .I(N__35908));
    LocalMux I__7218 (
            .O(N__35914),
            .I(N__35908));
    IoInMux I__7217 (
            .O(N__35913),
            .I(N__35905));
    Span4Mux_h I__7216 (
            .O(N__35908),
            .I(N__35901));
    LocalMux I__7215 (
            .O(N__35905),
            .I(N__35897));
    CEMux I__7214 (
            .O(N__35904),
            .I(N__35894));
    Span4Mux_v I__7213 (
            .O(N__35901),
            .I(N__35891));
    CEMux I__7212 (
            .O(N__35900),
            .I(N__35888));
    Span4Mux_s1_v I__7211 (
            .O(N__35897),
            .I(N__35885));
    LocalMux I__7210 (
            .O(N__35894),
            .I(N__35882));
    Span4Mux_v I__7209 (
            .O(N__35891),
            .I(N__35877));
    LocalMux I__7208 (
            .O(N__35888),
            .I(N__35877));
    Sp12to4 I__7207 (
            .O(N__35885),
            .I(N__35874));
    Span4Mux_v I__7206 (
            .O(N__35882),
            .I(N__35871));
    Span4Mux_h I__7205 (
            .O(N__35877),
            .I(N__35868));
    Span12Mux_h I__7204 (
            .O(N__35874),
            .I(N__35865));
    Span4Mux_v I__7203 (
            .O(N__35871),
            .I(N__35862));
    Span4Mux_v I__7202 (
            .O(N__35868),
            .I(N__35859));
    Span12Mux_v I__7201 (
            .O(N__35865),
            .I(N__35856));
    Span4Mux_v I__7200 (
            .O(N__35862),
            .I(N__35853));
    Span4Mux_v I__7199 (
            .O(N__35859),
            .I(N__35850));
    Odrv12 I__7198 (
            .O(N__35856),
            .I(red_c_i));
    Odrv4 I__7197 (
            .O(N__35853),
            .I(red_c_i));
    Odrv4 I__7196 (
            .O(N__35850),
            .I(red_c_i));
    InMux I__7195 (
            .O(N__35843),
            .I(N__35840));
    LocalMux I__7194 (
            .O(N__35840),
            .I(N__35837));
    Odrv4 I__7193 (
            .O(N__35837),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    CascadeMux I__7192 (
            .O(N__35834),
            .I(\phase_controller_inst2.start_timer_hc_RNO_0_0_cascade_ ));
    InMux I__7191 (
            .O(N__35831),
            .I(N__35828));
    LocalMux I__7190 (
            .O(N__35828),
            .I(N__35823));
    InMux I__7189 (
            .O(N__35827),
            .I(N__35819));
    InMux I__7188 (
            .O(N__35826),
            .I(N__35816));
    Span4Mux_v I__7187 (
            .O(N__35823),
            .I(N__35813));
    CascadeMux I__7186 (
            .O(N__35822),
            .I(N__35810));
    LocalMux I__7185 (
            .O(N__35819),
            .I(N__35805));
    LocalMux I__7184 (
            .O(N__35816),
            .I(N__35805));
    Span4Mux_v I__7183 (
            .O(N__35813),
            .I(N__35802));
    InMux I__7182 (
            .O(N__35810),
            .I(N__35799));
    Span4Mux_h I__7181 (
            .O(N__35805),
            .I(N__35796));
    Odrv4 I__7180 (
            .O(N__35802),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__7179 (
            .O(N__35799),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__7178 (
            .O(N__35796),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__7177 (
            .O(N__35789),
            .I(N__35786));
    LocalMux I__7176 (
            .O(N__35786),
            .I(N__35782));
    InMux I__7175 (
            .O(N__35785),
            .I(N__35778));
    Span4Mux_v I__7174 (
            .O(N__35782),
            .I(N__35775));
    InMux I__7173 (
            .O(N__35781),
            .I(N__35772));
    LocalMux I__7172 (
            .O(N__35778),
            .I(N__35765));
    Sp12to4 I__7171 (
            .O(N__35775),
            .I(N__35765));
    LocalMux I__7170 (
            .O(N__35772),
            .I(N__35765));
    Odrv12 I__7169 (
            .O(N__35765),
            .I(il_max_comp2_D2));
    InMux I__7168 (
            .O(N__35762),
            .I(N__35759));
    LocalMux I__7167 (
            .O(N__35759),
            .I(N__35756));
    Span4Mux_h I__7166 (
            .O(N__35756),
            .I(N__35753));
    Span4Mux_h I__7165 (
            .O(N__35753),
            .I(N__35749));
    CascadeMux I__7164 (
            .O(N__35752),
            .I(N__35746));
    Span4Mux_v I__7163 (
            .O(N__35749),
            .I(N__35742));
    InMux I__7162 (
            .O(N__35746),
            .I(N__35737));
    InMux I__7161 (
            .O(N__35745),
            .I(N__35737));
    Odrv4 I__7160 (
            .O(N__35742),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__7159 (
            .O(N__35737),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__7158 (
            .O(N__35732),
            .I(N__35729));
    LocalMux I__7157 (
            .O(N__35729),
            .I(N__35726));
    Odrv4 I__7156 (
            .O(N__35726),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__7155 (
            .O(N__35723),
            .I(N__35720));
    LocalMux I__7154 (
            .O(N__35720),
            .I(N__35716));
    InMux I__7153 (
            .O(N__35719),
            .I(N__35713));
    Odrv4 I__7152 (
            .O(N__35716),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__7151 (
            .O(N__35713),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__7150 (
            .O(N__35708),
            .I(\phase_controller_inst2.stoper_hc.time_passed11_cascade_ ));
    InMux I__7149 (
            .O(N__35705),
            .I(N__35702));
    LocalMux I__7148 (
            .O(N__35702),
            .I(N__35699));
    Span4Mux_h I__7147 (
            .O(N__35699),
            .I(N__35696));
    Odrv4 I__7146 (
            .O(N__35696),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__7145 (
            .O(N__35693),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__7144 (
            .O(N__35690),
            .I(N__35687));
    InMux I__7143 (
            .O(N__35687),
            .I(N__35684));
    LocalMux I__7142 (
            .O(N__35684),
            .I(N__35680));
    InMux I__7141 (
            .O(N__35683),
            .I(N__35676));
    Span4Mux_v I__7140 (
            .O(N__35680),
            .I(N__35673));
    InMux I__7139 (
            .O(N__35679),
            .I(N__35670));
    LocalMux I__7138 (
            .O(N__35676),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7137 (
            .O(N__35673),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__7136 (
            .O(N__35670),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__7135 (
            .O(N__35663),
            .I(N__35660));
    LocalMux I__7134 (
            .O(N__35660),
            .I(N__35657));
    Span4Mux_h I__7133 (
            .O(N__35657),
            .I(N__35654));
    Odrv4 I__7132 (
            .O(N__35654),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__7131 (
            .O(N__35651),
            .I(N__35648));
    LocalMux I__7130 (
            .O(N__35648),
            .I(N__35645));
    Span4Mux_h I__7129 (
            .O(N__35645),
            .I(N__35641));
    InMux I__7128 (
            .O(N__35644),
            .I(N__35638));
    Odrv4 I__7127 (
            .O(N__35641),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__7126 (
            .O(N__35638),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__7125 (
            .O(N__35633),
            .I(N__35626));
    InMux I__7124 (
            .O(N__35632),
            .I(N__35626));
    InMux I__7123 (
            .O(N__35631),
            .I(N__35623));
    LocalMux I__7122 (
            .O(N__35626),
            .I(N__35620));
    LocalMux I__7121 (
            .O(N__35623),
            .I(N__35616));
    Span4Mux_v I__7120 (
            .O(N__35620),
            .I(N__35613));
    InMux I__7119 (
            .O(N__35619),
            .I(N__35610));
    Span4Mux_v I__7118 (
            .O(N__35616),
            .I(N__35602));
    Span4Mux_h I__7117 (
            .O(N__35613),
            .I(N__35602));
    LocalMux I__7116 (
            .O(N__35610),
            .I(N__35602));
    InMux I__7115 (
            .O(N__35609),
            .I(N__35598));
    Span4Mux_h I__7114 (
            .O(N__35602),
            .I(N__35595));
    InMux I__7113 (
            .O(N__35601),
            .I(N__35592));
    LocalMux I__7112 (
            .O(N__35598),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__7111 (
            .O(N__35595),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__7110 (
            .O(N__35592),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__7109 (
            .O(N__35585),
            .I(N__35575));
    CascadeMux I__7108 (
            .O(N__35584),
            .I(N__35568));
    CascadeMux I__7107 (
            .O(N__35583),
            .I(N__35565));
    CascadeMux I__7106 (
            .O(N__35582),
            .I(N__35562));
    CascadeMux I__7105 (
            .O(N__35581),
            .I(N__35559));
    CascadeMux I__7104 (
            .O(N__35580),
            .I(N__35556));
    CascadeMux I__7103 (
            .O(N__35579),
            .I(N__35553));
    CascadeMux I__7102 (
            .O(N__35578),
            .I(N__35550));
    InMux I__7101 (
            .O(N__35575),
            .I(N__35537));
    InMux I__7100 (
            .O(N__35574),
            .I(N__35537));
    CascadeMux I__7099 (
            .O(N__35573),
            .I(N__35534));
    CascadeMux I__7098 (
            .O(N__35572),
            .I(N__35531));
    CascadeMux I__7097 (
            .O(N__35571),
            .I(N__35528));
    InMux I__7096 (
            .O(N__35568),
            .I(N__35520));
    InMux I__7095 (
            .O(N__35565),
            .I(N__35520));
    InMux I__7094 (
            .O(N__35562),
            .I(N__35520));
    InMux I__7093 (
            .O(N__35559),
            .I(N__35503));
    InMux I__7092 (
            .O(N__35556),
            .I(N__35503));
    InMux I__7091 (
            .O(N__35553),
            .I(N__35503));
    InMux I__7090 (
            .O(N__35550),
            .I(N__35503));
    InMux I__7089 (
            .O(N__35549),
            .I(N__35503));
    InMux I__7088 (
            .O(N__35548),
            .I(N__35503));
    InMux I__7087 (
            .O(N__35547),
            .I(N__35503));
    InMux I__7086 (
            .O(N__35546),
            .I(N__35503));
    InMux I__7085 (
            .O(N__35545),
            .I(N__35493));
    InMux I__7084 (
            .O(N__35544),
            .I(N__35493));
    InMux I__7083 (
            .O(N__35543),
            .I(N__35493));
    InMux I__7082 (
            .O(N__35542),
            .I(N__35493));
    LocalMux I__7081 (
            .O(N__35537),
            .I(N__35488));
    InMux I__7080 (
            .O(N__35534),
            .I(N__35479));
    InMux I__7079 (
            .O(N__35531),
            .I(N__35479));
    InMux I__7078 (
            .O(N__35528),
            .I(N__35479));
    InMux I__7077 (
            .O(N__35527),
            .I(N__35479));
    LocalMux I__7076 (
            .O(N__35520),
            .I(N__35474));
    LocalMux I__7075 (
            .O(N__35503),
            .I(N__35474));
    InMux I__7074 (
            .O(N__35502),
            .I(N__35471));
    LocalMux I__7073 (
            .O(N__35493),
            .I(N__35468));
    InMux I__7072 (
            .O(N__35492),
            .I(N__35463));
    InMux I__7071 (
            .O(N__35491),
            .I(N__35463));
    Span4Mux_v I__7070 (
            .O(N__35488),
            .I(N__35460));
    LocalMux I__7069 (
            .O(N__35479),
            .I(N__35455));
    Span4Mux_v I__7068 (
            .O(N__35474),
            .I(N__35455));
    LocalMux I__7067 (
            .O(N__35471),
            .I(N__35450));
    Span4Mux_h I__7066 (
            .O(N__35468),
            .I(N__35450));
    LocalMux I__7065 (
            .O(N__35463),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7064 (
            .O(N__35460),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7063 (
            .O(N__35455),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7062 (
            .O(N__35450),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__7061 (
            .O(N__35441),
            .I(N__35407));
    InMux I__7060 (
            .O(N__35440),
            .I(N__35407));
    InMux I__7059 (
            .O(N__35439),
            .I(N__35407));
    InMux I__7058 (
            .O(N__35438),
            .I(N__35407));
    InMux I__7057 (
            .O(N__35437),
            .I(N__35407));
    InMux I__7056 (
            .O(N__35436),
            .I(N__35407));
    InMux I__7055 (
            .O(N__35435),
            .I(N__35407));
    InMux I__7054 (
            .O(N__35434),
            .I(N__35390));
    InMux I__7053 (
            .O(N__35433),
            .I(N__35390));
    InMux I__7052 (
            .O(N__35432),
            .I(N__35390));
    InMux I__7051 (
            .O(N__35431),
            .I(N__35390));
    InMux I__7050 (
            .O(N__35430),
            .I(N__35390));
    InMux I__7049 (
            .O(N__35429),
            .I(N__35390));
    InMux I__7048 (
            .O(N__35428),
            .I(N__35390));
    InMux I__7047 (
            .O(N__35427),
            .I(N__35390));
    InMux I__7046 (
            .O(N__35426),
            .I(N__35381));
    InMux I__7045 (
            .O(N__35425),
            .I(N__35381));
    InMux I__7044 (
            .O(N__35424),
            .I(N__35381));
    InMux I__7043 (
            .O(N__35423),
            .I(N__35381));
    CascadeMux I__7042 (
            .O(N__35422),
            .I(N__35378));
    LocalMux I__7041 (
            .O(N__35407),
            .I(N__35368));
    LocalMux I__7040 (
            .O(N__35390),
            .I(N__35368));
    LocalMux I__7039 (
            .O(N__35381),
            .I(N__35368));
    InMux I__7038 (
            .O(N__35378),
            .I(N__35365));
    InMux I__7037 (
            .O(N__35377),
            .I(N__35362));
    InMux I__7036 (
            .O(N__35376),
            .I(N__35359));
    CascadeMux I__7035 (
            .O(N__35375),
            .I(N__35356));
    Span4Mux_v I__7034 (
            .O(N__35368),
            .I(N__35352));
    LocalMux I__7033 (
            .O(N__35365),
            .I(N__35345));
    LocalMux I__7032 (
            .O(N__35362),
            .I(N__35345));
    LocalMux I__7031 (
            .O(N__35359),
            .I(N__35345));
    InMux I__7030 (
            .O(N__35356),
            .I(N__35340));
    InMux I__7029 (
            .O(N__35355),
            .I(N__35340));
    Sp12to4 I__7028 (
            .O(N__35352),
            .I(N__35335));
    Span12Mux_v I__7027 (
            .O(N__35345),
            .I(N__35335));
    LocalMux I__7026 (
            .O(N__35340),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__7025 (
            .O(N__35335),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__7024 (
            .O(N__35330),
            .I(N__35321));
    CascadeMux I__7023 (
            .O(N__35329),
            .I(N__35318));
    CascadeMux I__7022 (
            .O(N__35328),
            .I(N__35315));
    CascadeMux I__7021 (
            .O(N__35327),
            .I(N__35312));
    CascadeMux I__7020 (
            .O(N__35326),
            .I(N__35298));
    CascadeMux I__7019 (
            .O(N__35325),
            .I(N__35295));
    CascadeMux I__7018 (
            .O(N__35324),
            .I(N__35292));
    InMux I__7017 (
            .O(N__35321),
            .I(N__35279));
    InMux I__7016 (
            .O(N__35318),
            .I(N__35279));
    InMux I__7015 (
            .O(N__35315),
            .I(N__35279));
    InMux I__7014 (
            .O(N__35312),
            .I(N__35279));
    InMux I__7013 (
            .O(N__35311),
            .I(N__35270));
    InMux I__7012 (
            .O(N__35310),
            .I(N__35270));
    InMux I__7011 (
            .O(N__35309),
            .I(N__35270));
    InMux I__7010 (
            .O(N__35308),
            .I(N__35270));
    InMux I__7009 (
            .O(N__35307),
            .I(N__35255));
    InMux I__7008 (
            .O(N__35306),
            .I(N__35255));
    InMux I__7007 (
            .O(N__35305),
            .I(N__35255));
    InMux I__7006 (
            .O(N__35304),
            .I(N__35255));
    InMux I__7005 (
            .O(N__35303),
            .I(N__35255));
    InMux I__7004 (
            .O(N__35302),
            .I(N__35255));
    InMux I__7003 (
            .O(N__35301),
            .I(N__35255));
    InMux I__7002 (
            .O(N__35298),
            .I(N__35250));
    InMux I__7001 (
            .O(N__35295),
            .I(N__35250));
    InMux I__7000 (
            .O(N__35292),
            .I(N__35245));
    InMux I__6999 (
            .O(N__35291),
            .I(N__35245));
    InMux I__6998 (
            .O(N__35290),
            .I(N__35242));
    InMux I__6997 (
            .O(N__35289),
            .I(N__35239));
    InMux I__6996 (
            .O(N__35288),
            .I(N__35236));
    LocalMux I__6995 (
            .O(N__35279),
            .I(N__35229));
    LocalMux I__6994 (
            .O(N__35270),
            .I(N__35229));
    LocalMux I__6993 (
            .O(N__35255),
            .I(N__35229));
    LocalMux I__6992 (
            .O(N__35250),
            .I(N__35226));
    LocalMux I__6991 (
            .O(N__35245),
            .I(N__35223));
    LocalMux I__6990 (
            .O(N__35242),
            .I(N__35216));
    LocalMux I__6989 (
            .O(N__35239),
            .I(N__35216));
    LocalMux I__6988 (
            .O(N__35236),
            .I(N__35216));
    Span4Mux_v I__6987 (
            .O(N__35229),
            .I(N__35211));
    Span4Mux_h I__6986 (
            .O(N__35226),
            .I(N__35206));
    Span4Mux_h I__6985 (
            .O(N__35223),
            .I(N__35206));
    Span4Mux_v I__6984 (
            .O(N__35216),
            .I(N__35203));
    InMux I__6983 (
            .O(N__35215),
            .I(N__35198));
    InMux I__6982 (
            .O(N__35214),
            .I(N__35198));
    Span4Mux_h I__6981 (
            .O(N__35211),
            .I(N__35195));
    Span4Mux_h I__6980 (
            .O(N__35206),
            .I(N__35192));
    Span4Mux_h I__6979 (
            .O(N__35203),
            .I(N__35189));
    LocalMux I__6978 (
            .O(N__35198),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6977 (
            .O(N__35195),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6976 (
            .O(N__35192),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6975 (
            .O(N__35189),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__6974 (
            .O(N__35180),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__6973 (
            .O(N__35177),
            .I(N__35174));
    InMux I__6972 (
            .O(N__35174),
            .I(N__35171));
    LocalMux I__6971 (
            .O(N__35171),
            .I(N__35166));
    CascadeMux I__6970 (
            .O(N__35170),
            .I(N__35163));
    InMux I__6969 (
            .O(N__35169),
            .I(N__35160));
    Span4Mux_v I__6968 (
            .O(N__35166),
            .I(N__35157));
    InMux I__6967 (
            .O(N__35163),
            .I(N__35154));
    LocalMux I__6966 (
            .O(N__35160),
            .I(N__35151));
    Odrv4 I__6965 (
            .O(N__35157),
            .I(measured_delay_tr_3));
    LocalMux I__6964 (
            .O(N__35154),
            .I(measured_delay_tr_3));
    Odrv4 I__6963 (
            .O(N__35151),
            .I(measured_delay_tr_3));
    InMux I__6962 (
            .O(N__35144),
            .I(N__35141));
    LocalMux I__6961 (
            .O(N__35141),
            .I(N__35137));
    InMux I__6960 (
            .O(N__35140),
            .I(N__35134));
    Span4Mux_v I__6959 (
            .O(N__35137),
            .I(N__35128));
    LocalMux I__6958 (
            .O(N__35134),
            .I(N__35128));
    InMux I__6957 (
            .O(N__35133),
            .I(N__35125));
    Odrv4 I__6956 (
            .O(N__35128),
            .I(\phase_controller_inst1.stoper_tr.N_248 ));
    LocalMux I__6955 (
            .O(N__35125),
            .I(\phase_controller_inst1.stoper_tr.N_248 ));
    CascadeMux I__6954 (
            .O(N__35120),
            .I(N__35117));
    InMux I__6953 (
            .O(N__35117),
            .I(N__35114));
    LocalMux I__6952 (
            .O(N__35114),
            .I(N__35110));
    CascadeMux I__6951 (
            .O(N__35113),
            .I(N__35107));
    Span4Mux_v I__6950 (
            .O(N__35110),
            .I(N__35104));
    InMux I__6949 (
            .O(N__35107),
            .I(N__35101));
    Odrv4 I__6948 (
            .O(N__35104),
            .I(measured_delay_tr_1));
    LocalMux I__6947 (
            .O(N__35101),
            .I(measured_delay_tr_1));
    InMux I__6946 (
            .O(N__35096),
            .I(N__35093));
    LocalMux I__6945 (
            .O(N__35093),
            .I(N__35089));
    InMux I__6944 (
            .O(N__35092),
            .I(N__35086));
    Span4Mux_v I__6943 (
            .O(N__35089),
            .I(N__35082));
    LocalMux I__6942 (
            .O(N__35086),
            .I(N__35079));
    InMux I__6941 (
            .O(N__35085),
            .I(N__35076));
    Odrv4 I__6940 (
            .O(N__35082),
            .I(measured_delay_tr_11));
    Odrv4 I__6939 (
            .O(N__35079),
            .I(measured_delay_tr_11));
    LocalMux I__6938 (
            .O(N__35076),
            .I(measured_delay_tr_11));
    InMux I__6937 (
            .O(N__35069),
            .I(N__35066));
    LocalMux I__6936 (
            .O(N__35066),
            .I(N__35061));
    InMux I__6935 (
            .O(N__35065),
            .I(N__35058));
    InMux I__6934 (
            .O(N__35064),
            .I(N__35055));
    Span4Mux_v I__6933 (
            .O(N__35061),
            .I(N__35052));
    LocalMux I__6932 (
            .O(N__35058),
            .I(N__35049));
    LocalMux I__6931 (
            .O(N__35055),
            .I(N__35046));
    Odrv4 I__6930 (
            .O(N__35052),
            .I(measured_delay_tr_9));
    Odrv4 I__6929 (
            .O(N__35049),
            .I(measured_delay_tr_9));
    Odrv4 I__6928 (
            .O(N__35046),
            .I(measured_delay_tr_9));
    InMux I__6927 (
            .O(N__35039),
            .I(N__35034));
    InMux I__6926 (
            .O(N__35038),
            .I(N__35030));
    InMux I__6925 (
            .O(N__35037),
            .I(N__35027));
    LocalMux I__6924 (
            .O(N__35034),
            .I(N__35024));
    InMux I__6923 (
            .O(N__35033),
            .I(N__35021));
    LocalMux I__6922 (
            .O(N__35030),
            .I(N__35016));
    LocalMux I__6921 (
            .O(N__35027),
            .I(N__35016));
    Odrv4 I__6920 (
            .O(N__35024),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    LocalMux I__6919 (
            .O(N__35021),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    Odrv12 I__6918 (
            .O(N__35016),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    InMux I__6917 (
            .O(N__35009),
            .I(N__35005));
    InMux I__6916 (
            .O(N__35008),
            .I(N__35002));
    LocalMux I__6915 (
            .O(N__35005),
            .I(N__34999));
    LocalMux I__6914 (
            .O(N__35002),
            .I(N__34995));
    Span12Mux_v I__6913 (
            .O(N__34999),
            .I(N__34992));
    InMux I__6912 (
            .O(N__34998),
            .I(N__34989));
    Odrv4 I__6911 (
            .O(N__34995),
            .I(measured_delay_tr_6));
    Odrv12 I__6910 (
            .O(N__34992),
            .I(measured_delay_tr_6));
    LocalMux I__6909 (
            .O(N__34989),
            .I(measured_delay_tr_6));
    InMux I__6908 (
            .O(N__34982),
            .I(N__34979));
    LocalMux I__6907 (
            .O(N__34979),
            .I(N__34975));
    InMux I__6906 (
            .O(N__34978),
            .I(N__34972));
    Span4Mux_v I__6905 (
            .O(N__34975),
            .I(N__34966));
    LocalMux I__6904 (
            .O(N__34972),
            .I(N__34966));
    InMux I__6903 (
            .O(N__34971),
            .I(N__34963));
    Span4Mux_v I__6902 (
            .O(N__34966),
            .I(N__34960));
    LocalMux I__6901 (
            .O(N__34963),
            .I(N__34957));
    Odrv4 I__6900 (
            .O(N__34960),
            .I(measured_delay_tr_2));
    Odrv4 I__6899 (
            .O(N__34957),
            .I(measured_delay_tr_2));
    InMux I__6898 (
            .O(N__34952),
            .I(N__34948));
    InMux I__6897 (
            .O(N__34951),
            .I(N__34945));
    LocalMux I__6896 (
            .O(N__34948),
            .I(N__34940));
    LocalMux I__6895 (
            .O(N__34945),
            .I(N__34940));
    Span4Mux_v I__6894 (
            .O(N__34940),
            .I(N__34935));
    InMux I__6893 (
            .O(N__34939),
            .I(N__34932));
    InMux I__6892 (
            .O(N__34938),
            .I(N__34929));
    Odrv4 I__6891 (
            .O(N__34935),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    LocalMux I__6890 (
            .O(N__34932),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    LocalMux I__6889 (
            .O(N__34929),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    InMux I__6888 (
            .O(N__34922),
            .I(N__34919));
    LocalMux I__6887 (
            .O(N__34919),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ));
    InMux I__6886 (
            .O(N__34916),
            .I(N__34913));
    LocalMux I__6885 (
            .O(N__34913),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ));
    InMux I__6884 (
            .O(N__34910),
            .I(N__34907));
    LocalMux I__6883 (
            .O(N__34907),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ));
    CascadeMux I__6882 (
            .O(N__34904),
            .I(N__34901));
    InMux I__6881 (
            .O(N__34901),
            .I(N__34898));
    LocalMux I__6880 (
            .O(N__34898),
            .I(N__34895));
    Odrv12 I__6879 (
            .O(N__34895),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__6878 (
            .O(N__34892),
            .I(N__34889));
    LocalMux I__6877 (
            .O(N__34889),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ));
    InMux I__6876 (
            .O(N__34886),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__6875 (
            .O(N__34883),
            .I(N__34880));
    InMux I__6874 (
            .O(N__34880),
            .I(N__34877));
    LocalMux I__6873 (
            .O(N__34877),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__6872 (
            .O(N__34874),
            .I(N__34871));
    InMux I__6871 (
            .O(N__34871),
            .I(N__34868));
    LocalMux I__6870 (
            .O(N__34868),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__6869 (
            .O(N__34865),
            .I(N__34861));
    InMux I__6868 (
            .O(N__34864),
            .I(N__34857));
    LocalMux I__6867 (
            .O(N__34861),
            .I(N__34854));
    InMux I__6866 (
            .O(N__34860),
            .I(N__34851));
    LocalMux I__6865 (
            .O(N__34857),
            .I(N__34848));
    Odrv4 I__6864 (
            .O(N__34854),
            .I(measured_delay_tr_5));
    LocalMux I__6863 (
            .O(N__34851),
            .I(measured_delay_tr_5));
    Odrv4 I__6862 (
            .O(N__34848),
            .I(measured_delay_tr_5));
    CascadeMux I__6861 (
            .O(N__34841),
            .I(N__34838));
    InMux I__6860 (
            .O(N__34838),
            .I(N__34835));
    LocalMux I__6859 (
            .O(N__34835),
            .I(N__34832));
    Odrv12 I__6858 (
            .O(N__34832),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    InMux I__6857 (
            .O(N__34829),
            .I(N__34826));
    LocalMux I__6856 (
            .O(N__34826),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__6855 (
            .O(N__34823),
            .I(N__34820));
    InMux I__6854 (
            .O(N__34820),
            .I(N__34817));
    LocalMux I__6853 (
            .O(N__34817),
            .I(N__34814));
    Odrv4 I__6852 (
            .O(N__34814),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__6851 (
            .O(N__34811),
            .I(N__34808));
    LocalMux I__6850 (
            .O(N__34808),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__6849 (
            .O(N__34805),
            .I(N__34802));
    LocalMux I__6848 (
            .O(N__34802),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__6847 (
            .O(N__34799),
            .I(N__34796));
    InMux I__6846 (
            .O(N__34796),
            .I(N__34793));
    LocalMux I__6845 (
            .O(N__34793),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__6844 (
            .O(N__34790),
            .I(N__34787));
    LocalMux I__6843 (
            .O(N__34787),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__6842 (
            .O(N__34784),
            .I(N__34781));
    InMux I__6841 (
            .O(N__34781),
            .I(N__34778));
    LocalMux I__6840 (
            .O(N__34778),
            .I(N__34775));
    Span4Mux_h I__6839 (
            .O(N__34775),
            .I(N__34772));
    Odrv4 I__6838 (
            .O(N__34772),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__6837 (
            .O(N__34769),
            .I(N__34766));
    LocalMux I__6836 (
            .O(N__34766),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__6835 (
            .O(N__34763),
            .I(N__34760));
    LocalMux I__6834 (
            .O(N__34760),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__6833 (
            .O(N__34757),
            .I(N__34754));
    LocalMux I__6832 (
            .O(N__34754),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__6831 (
            .O(N__34751),
            .I(N__34748));
    InMux I__6830 (
            .O(N__34748),
            .I(N__34745));
    LocalMux I__6829 (
            .O(N__34745),
            .I(N__34742));
    Span4Mux_v I__6828 (
            .O(N__34742),
            .I(N__34739));
    Odrv4 I__6827 (
            .O(N__34739),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    InMux I__6826 (
            .O(N__34736),
            .I(N__34733));
    LocalMux I__6825 (
            .O(N__34733),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__6824 (
            .O(N__34730),
            .I(N__34727));
    LocalMux I__6823 (
            .O(N__34727),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__6822 (
            .O(N__34724),
            .I(N__34721));
    InMux I__6821 (
            .O(N__34721),
            .I(N__34718));
    LocalMux I__6820 (
            .O(N__34718),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__6819 (
            .O(N__34715),
            .I(N__34712));
    InMux I__6818 (
            .O(N__34712),
            .I(N__34709));
    LocalMux I__6817 (
            .O(N__34709),
            .I(N__34706));
    Odrv4 I__6816 (
            .O(N__34706),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    InMux I__6815 (
            .O(N__34703),
            .I(N__34700));
    LocalMux I__6814 (
            .O(N__34700),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__6813 (
            .O(N__34697),
            .I(N__34694));
    InMux I__6812 (
            .O(N__34694),
            .I(N__34691));
    LocalMux I__6811 (
            .O(N__34691),
            .I(N__34688));
    Odrv12 I__6810 (
            .O(N__34688),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__6809 (
            .O(N__34685),
            .I(N__34682));
    LocalMux I__6808 (
            .O(N__34682),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__6807 (
            .O(N__34679),
            .I(N__34676));
    LocalMux I__6806 (
            .O(N__34676),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__6805 (
            .O(N__34673),
            .I(N__34670));
    LocalMux I__6804 (
            .O(N__34670),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__6803 (
            .O(N__34667),
            .I(N__34664));
    InMux I__6802 (
            .O(N__34664),
            .I(N__34661));
    LocalMux I__6801 (
            .O(N__34661),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__6800 (
            .O(N__34658),
            .I(N__34655));
    InMux I__6799 (
            .O(N__34655),
            .I(N__34652));
    LocalMux I__6798 (
            .O(N__34652),
            .I(N__34649));
    Span4Mux_h I__6797 (
            .O(N__34649),
            .I(N__34646));
    Odrv4 I__6796 (
            .O(N__34646),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    InMux I__6795 (
            .O(N__34643),
            .I(N__34640));
    LocalMux I__6794 (
            .O(N__34640),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__6793 (
            .O(N__34637),
            .I(N__34634));
    InMux I__6792 (
            .O(N__34634),
            .I(N__34631));
    LocalMux I__6791 (
            .O(N__34631),
            .I(N__34628));
    Span4Mux_h I__6790 (
            .O(N__34628),
            .I(N__34625));
    Odrv4 I__6789 (
            .O(N__34625),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__6788 (
            .O(N__34622),
            .I(N__34619));
    LocalMux I__6787 (
            .O(N__34619),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__6786 (
            .O(N__34616),
            .I(N__34613));
    InMux I__6785 (
            .O(N__34613),
            .I(N__34603));
    InMux I__6784 (
            .O(N__34612),
            .I(N__34603));
    CascadeMux I__6783 (
            .O(N__34611),
            .I(N__34600));
    InMux I__6782 (
            .O(N__34610),
            .I(N__34593));
    InMux I__6781 (
            .O(N__34609),
            .I(N__34593));
    InMux I__6780 (
            .O(N__34608),
            .I(N__34593));
    LocalMux I__6779 (
            .O(N__34603),
            .I(N__34590));
    InMux I__6778 (
            .O(N__34600),
            .I(N__34587));
    LocalMux I__6777 (
            .O(N__34593),
            .I(N__34584));
    Span4Mux_h I__6776 (
            .O(N__34590),
            .I(N__34581));
    LocalMux I__6775 (
            .O(N__34587),
            .I(state_3));
    Odrv12 I__6774 (
            .O(N__34584),
            .I(state_3));
    Odrv4 I__6773 (
            .O(N__34581),
            .I(state_3));
    IoInMux I__6772 (
            .O(N__34574),
            .I(N__34571));
    LocalMux I__6771 (
            .O(N__34571),
            .I(N__34568));
    Span4Mux_s1_v I__6770 (
            .O(N__34568),
            .I(N__34564));
    CascadeMux I__6769 (
            .O(N__34567),
            .I(N__34561));
    Span4Mux_v I__6768 (
            .O(N__34564),
            .I(N__34557));
    InMux I__6767 (
            .O(N__34561),
            .I(N__34552));
    InMux I__6766 (
            .O(N__34560),
            .I(N__34552));
    Odrv4 I__6765 (
            .O(N__34557),
            .I(s1_phy_c));
    LocalMux I__6764 (
            .O(N__34552),
            .I(s1_phy_c));
    InMux I__6763 (
            .O(N__34547),
            .I(N__34537));
    InMux I__6762 (
            .O(N__34546),
            .I(N__34537));
    InMux I__6761 (
            .O(N__34545),
            .I(N__34537));
    InMux I__6760 (
            .O(N__34544),
            .I(N__34534));
    LocalMux I__6759 (
            .O(N__34537),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6758 (
            .O(N__34534),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    IoInMux I__6757 (
            .O(N__34529),
            .I(N__34526));
    LocalMux I__6756 (
            .O(N__34526),
            .I(N__34523));
    Odrv12 I__6755 (
            .O(N__34523),
            .I(\current_shift_inst.timer_s1.N_181_i ));
    IoInMux I__6754 (
            .O(N__34520),
            .I(N__34517));
    LocalMux I__6753 (
            .O(N__34517),
            .I(N__34514));
    Odrv12 I__6752 (
            .O(N__34514),
            .I(s2_phy_c));
    CascadeMux I__6751 (
            .O(N__34511),
            .I(\phase_controller_inst2.stoper_tr.time_passed11_cascade_ ));
    CascadeMux I__6750 (
            .O(N__34508),
            .I(N__34503));
    InMux I__6749 (
            .O(N__34507),
            .I(N__34499));
    CascadeMux I__6748 (
            .O(N__34506),
            .I(N__34496));
    InMux I__6747 (
            .O(N__34503),
            .I(N__34493));
    CascadeMux I__6746 (
            .O(N__34502),
            .I(N__34490));
    LocalMux I__6745 (
            .O(N__34499),
            .I(N__34487));
    InMux I__6744 (
            .O(N__34496),
            .I(N__34484));
    LocalMux I__6743 (
            .O(N__34493),
            .I(N__34481));
    InMux I__6742 (
            .O(N__34490),
            .I(N__34478));
    Span4Mux_h I__6741 (
            .O(N__34487),
            .I(N__34475));
    LocalMux I__6740 (
            .O(N__34484),
            .I(N__34472));
    Span4Mux_h I__6739 (
            .O(N__34481),
            .I(N__34467));
    LocalMux I__6738 (
            .O(N__34478),
            .I(N__34467));
    Span4Mux_v I__6737 (
            .O(N__34475),
            .I(N__34463));
    Span4Mux_h I__6736 (
            .O(N__34472),
            .I(N__34458));
    Span4Mux_h I__6735 (
            .O(N__34467),
            .I(N__34458));
    InMux I__6734 (
            .O(N__34466),
            .I(N__34455));
    Span4Mux_h I__6733 (
            .O(N__34463),
            .I(N__34452));
    Span4Mux_v I__6732 (
            .O(N__34458),
            .I(N__34449));
    LocalMux I__6731 (
            .O(N__34455),
            .I(measured_delay_hc_13));
    Odrv4 I__6730 (
            .O(N__34452),
            .I(measured_delay_hc_13));
    Odrv4 I__6729 (
            .O(N__34449),
            .I(measured_delay_hc_13));
    CascadeMux I__6728 (
            .O(N__34442),
            .I(N__34439));
    InMux I__6727 (
            .O(N__34439),
            .I(N__34436));
    LocalMux I__6726 (
            .O(N__34436),
            .I(N__34433));
    Odrv12 I__6725 (
            .O(N__34433),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__6724 (
            .O(N__34430),
            .I(N__34425));
    InMux I__6723 (
            .O(N__34429),
            .I(N__34421));
    InMux I__6722 (
            .O(N__34428),
            .I(N__34418));
    LocalMux I__6721 (
            .O(N__34425),
            .I(N__34415));
    InMux I__6720 (
            .O(N__34424),
            .I(N__34412));
    LocalMux I__6719 (
            .O(N__34421),
            .I(N__34409));
    LocalMux I__6718 (
            .O(N__34418),
            .I(N__34406));
    Span4Mux_h I__6717 (
            .O(N__34415),
            .I(N__34401));
    LocalMux I__6716 (
            .O(N__34412),
            .I(N__34401));
    Span4Mux_h I__6715 (
            .O(N__34409),
            .I(N__34395));
    Span4Mux_h I__6714 (
            .O(N__34406),
            .I(N__34395));
    Span4Mux_h I__6713 (
            .O(N__34401),
            .I(N__34392));
    InMux I__6712 (
            .O(N__34400),
            .I(N__34389));
    Span4Mux_v I__6711 (
            .O(N__34395),
            .I(N__34386));
    Odrv4 I__6710 (
            .O(N__34392),
            .I(measured_delay_hc_15));
    LocalMux I__6709 (
            .O(N__34389),
            .I(measured_delay_hc_15));
    Odrv4 I__6708 (
            .O(N__34386),
            .I(measured_delay_hc_15));
    CascadeMux I__6707 (
            .O(N__34379),
            .I(N__34376));
    InMux I__6706 (
            .O(N__34376),
            .I(N__34373));
    LocalMux I__6705 (
            .O(N__34373),
            .I(N__34370));
    Span4Mux_v I__6704 (
            .O(N__34370),
            .I(N__34367));
    Odrv4 I__6703 (
            .O(N__34367),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__6702 (
            .O(N__34364),
            .I(N__34353));
    CascadeMux I__6701 (
            .O(N__34363),
            .I(N__34350));
    CascadeMux I__6700 (
            .O(N__34362),
            .I(N__34347));
    CascadeMux I__6699 (
            .O(N__34361),
            .I(N__34344));
    InMux I__6698 (
            .O(N__34360),
            .I(N__34329));
    InMux I__6697 (
            .O(N__34359),
            .I(N__34329));
    InMux I__6696 (
            .O(N__34358),
            .I(N__34329));
    InMux I__6695 (
            .O(N__34357),
            .I(N__34326));
    InMux I__6694 (
            .O(N__34356),
            .I(N__34309));
    InMux I__6693 (
            .O(N__34353),
            .I(N__34309));
    InMux I__6692 (
            .O(N__34350),
            .I(N__34309));
    InMux I__6691 (
            .O(N__34347),
            .I(N__34309));
    InMux I__6690 (
            .O(N__34344),
            .I(N__34309));
    InMux I__6689 (
            .O(N__34343),
            .I(N__34309));
    InMux I__6688 (
            .O(N__34342),
            .I(N__34309));
    InMux I__6687 (
            .O(N__34341),
            .I(N__34309));
    InMux I__6686 (
            .O(N__34340),
            .I(N__34304));
    InMux I__6685 (
            .O(N__34339),
            .I(N__34304));
    CascadeMux I__6684 (
            .O(N__34338),
            .I(N__34300));
    CascadeMux I__6683 (
            .O(N__34337),
            .I(N__34297));
    CascadeMux I__6682 (
            .O(N__34336),
            .I(N__34285));
    LocalMux I__6681 (
            .O(N__34329),
            .I(N__34277));
    LocalMux I__6680 (
            .O(N__34326),
            .I(N__34277));
    LocalMux I__6679 (
            .O(N__34309),
            .I(N__34277));
    LocalMux I__6678 (
            .O(N__34304),
            .I(N__34274));
    InMux I__6677 (
            .O(N__34303),
            .I(N__34271));
    InMux I__6676 (
            .O(N__34300),
            .I(N__34259));
    InMux I__6675 (
            .O(N__34297),
            .I(N__34259));
    InMux I__6674 (
            .O(N__34296),
            .I(N__34250));
    InMux I__6673 (
            .O(N__34295),
            .I(N__34250));
    InMux I__6672 (
            .O(N__34294),
            .I(N__34250));
    InMux I__6671 (
            .O(N__34293),
            .I(N__34250));
    InMux I__6670 (
            .O(N__34292),
            .I(N__34239));
    InMux I__6669 (
            .O(N__34291),
            .I(N__34239));
    InMux I__6668 (
            .O(N__34290),
            .I(N__34239));
    InMux I__6667 (
            .O(N__34289),
            .I(N__34239));
    InMux I__6666 (
            .O(N__34288),
            .I(N__34239));
    InMux I__6665 (
            .O(N__34285),
            .I(N__34234));
    InMux I__6664 (
            .O(N__34284),
            .I(N__34234));
    Span4Mux_v I__6663 (
            .O(N__34277),
            .I(N__34227));
    Span4Mux_v I__6662 (
            .O(N__34274),
            .I(N__34227));
    LocalMux I__6661 (
            .O(N__34271),
            .I(N__34227));
    InMux I__6660 (
            .O(N__34270),
            .I(N__34224));
    InMux I__6659 (
            .O(N__34269),
            .I(N__34211));
    InMux I__6658 (
            .O(N__34268),
            .I(N__34211));
    InMux I__6657 (
            .O(N__34267),
            .I(N__34211));
    InMux I__6656 (
            .O(N__34266),
            .I(N__34211));
    InMux I__6655 (
            .O(N__34265),
            .I(N__34211));
    InMux I__6654 (
            .O(N__34264),
            .I(N__34211));
    LocalMux I__6653 (
            .O(N__34259),
            .I(N__34206));
    LocalMux I__6652 (
            .O(N__34250),
            .I(N__34206));
    LocalMux I__6651 (
            .O(N__34239),
            .I(N__34203));
    LocalMux I__6650 (
            .O(N__34234),
            .I(N__34200));
    Span4Mux_h I__6649 (
            .O(N__34227),
            .I(N__34197));
    LocalMux I__6648 (
            .O(N__34224),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    LocalMux I__6647 (
            .O(N__34211),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    Odrv4 I__6646 (
            .O(N__34206),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    Odrv4 I__6645 (
            .O(N__34203),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    Odrv12 I__6644 (
            .O(N__34200),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    Odrv4 I__6643 (
            .O(N__34197),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    InMux I__6642 (
            .O(N__34184),
            .I(N__34178));
    InMux I__6641 (
            .O(N__34183),
            .I(N__34178));
    LocalMux I__6640 (
            .O(N__34178),
            .I(N__34162));
    InMux I__6639 (
            .O(N__34177),
            .I(N__34157));
    InMux I__6638 (
            .O(N__34176),
            .I(N__34157));
    InMux I__6637 (
            .O(N__34175),
            .I(N__34142));
    InMux I__6636 (
            .O(N__34174),
            .I(N__34142));
    InMux I__6635 (
            .O(N__34173),
            .I(N__34142));
    InMux I__6634 (
            .O(N__34172),
            .I(N__34142));
    InMux I__6633 (
            .O(N__34171),
            .I(N__34142));
    InMux I__6632 (
            .O(N__34170),
            .I(N__34142));
    InMux I__6631 (
            .O(N__34169),
            .I(N__34131));
    InMux I__6630 (
            .O(N__34168),
            .I(N__34131));
    InMux I__6629 (
            .O(N__34167),
            .I(N__34131));
    InMux I__6628 (
            .O(N__34166),
            .I(N__34131));
    InMux I__6627 (
            .O(N__34165),
            .I(N__34131));
    Span4Mux_h I__6626 (
            .O(N__34162),
            .I(N__34123));
    LocalMux I__6625 (
            .O(N__34157),
            .I(N__34123));
    InMux I__6624 (
            .O(N__34156),
            .I(N__34118));
    InMux I__6623 (
            .O(N__34155),
            .I(N__34118));
    LocalMux I__6622 (
            .O(N__34142),
            .I(N__34115));
    LocalMux I__6621 (
            .O(N__34131),
            .I(N__34112));
    InMux I__6620 (
            .O(N__34130),
            .I(N__34105));
    InMux I__6619 (
            .O(N__34129),
            .I(N__34105));
    InMux I__6618 (
            .O(N__34128),
            .I(N__34105));
    Span4Mux_h I__6617 (
            .O(N__34123),
            .I(N__34094));
    LocalMux I__6616 (
            .O(N__34118),
            .I(N__34091));
    Span4Mux_v I__6615 (
            .O(N__34115),
            .I(N__34084));
    Span4Mux_h I__6614 (
            .O(N__34112),
            .I(N__34084));
    LocalMux I__6613 (
            .O(N__34105),
            .I(N__34084));
    InMux I__6612 (
            .O(N__34104),
            .I(N__34067));
    InMux I__6611 (
            .O(N__34103),
            .I(N__34067));
    InMux I__6610 (
            .O(N__34102),
            .I(N__34067));
    InMux I__6609 (
            .O(N__34101),
            .I(N__34067));
    InMux I__6608 (
            .O(N__34100),
            .I(N__34067));
    InMux I__6607 (
            .O(N__34099),
            .I(N__34067));
    InMux I__6606 (
            .O(N__34098),
            .I(N__34067));
    InMux I__6605 (
            .O(N__34097),
            .I(N__34067));
    Odrv4 I__6604 (
            .O(N__34094),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt30 ));
    Odrv4 I__6603 (
            .O(N__34091),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt30 ));
    Odrv4 I__6602 (
            .O(N__34084),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt30 ));
    LocalMux I__6601 (
            .O(N__34067),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt30 ));
    CascadeMux I__6600 (
            .O(N__34058),
            .I(N__34055));
    InMux I__6599 (
            .O(N__34055),
            .I(N__34051));
    CascadeMux I__6598 (
            .O(N__34054),
            .I(N__34048));
    LocalMux I__6597 (
            .O(N__34051),
            .I(N__34045));
    InMux I__6596 (
            .O(N__34048),
            .I(N__34040));
    Span4Mux_v I__6595 (
            .O(N__34045),
            .I(N__34036));
    InMux I__6594 (
            .O(N__34044),
            .I(N__34031));
    InMux I__6593 (
            .O(N__34043),
            .I(N__34031));
    LocalMux I__6592 (
            .O(N__34040),
            .I(N__34028));
    InMux I__6591 (
            .O(N__34039),
            .I(N__34025));
    Span4Mux_h I__6590 (
            .O(N__34036),
            .I(N__34020));
    LocalMux I__6589 (
            .O(N__34031),
            .I(N__34020));
    Odrv4 I__6588 (
            .O(N__34028),
            .I(measured_delay_hc_2));
    LocalMux I__6587 (
            .O(N__34025),
            .I(measured_delay_hc_2));
    Odrv4 I__6586 (
            .O(N__34020),
            .I(measured_delay_hc_2));
    CascadeMux I__6585 (
            .O(N__34013),
            .I(N__34005));
    CascadeMux I__6584 (
            .O(N__34012),
            .I(N__33999));
    CascadeMux I__6583 (
            .O(N__34011),
            .I(N__33996));
    CascadeMux I__6582 (
            .O(N__34010),
            .I(N__33993));
    InMux I__6581 (
            .O(N__34009),
            .I(N__33987));
    InMux I__6580 (
            .O(N__34008),
            .I(N__33987));
    InMux I__6579 (
            .O(N__34005),
            .I(N__33976));
    InMux I__6578 (
            .O(N__34004),
            .I(N__33976));
    InMux I__6577 (
            .O(N__34003),
            .I(N__33976));
    InMux I__6576 (
            .O(N__34002),
            .I(N__33976));
    InMux I__6575 (
            .O(N__33999),
            .I(N__33967));
    InMux I__6574 (
            .O(N__33996),
            .I(N__33967));
    InMux I__6573 (
            .O(N__33993),
            .I(N__33967));
    InMux I__6572 (
            .O(N__33992),
            .I(N__33967));
    LocalMux I__6571 (
            .O(N__33987),
            .I(N__33964));
    CascadeMux I__6570 (
            .O(N__33986),
            .I(N__33952));
    CascadeMux I__6569 (
            .O(N__33985),
            .I(N__33949));
    LocalMux I__6568 (
            .O(N__33976),
            .I(N__33942));
    LocalMux I__6567 (
            .O(N__33967),
            .I(N__33937));
    Span4Mux_h I__6566 (
            .O(N__33964),
            .I(N__33937));
    CascadeMux I__6565 (
            .O(N__33963),
            .I(N__33932));
    CascadeMux I__6564 (
            .O(N__33962),
            .I(N__33929));
    CascadeMux I__6563 (
            .O(N__33961),
            .I(N__33924));
    CascadeMux I__6562 (
            .O(N__33960),
            .I(N__33918));
    CascadeMux I__6561 (
            .O(N__33959),
            .I(N__33915));
    CascadeMux I__6560 (
            .O(N__33958),
            .I(N__33912));
    InMux I__6559 (
            .O(N__33957),
            .I(N__33904));
    InMux I__6558 (
            .O(N__33956),
            .I(N__33887));
    InMux I__6557 (
            .O(N__33955),
            .I(N__33887));
    InMux I__6556 (
            .O(N__33952),
            .I(N__33887));
    InMux I__6555 (
            .O(N__33949),
            .I(N__33887));
    InMux I__6554 (
            .O(N__33948),
            .I(N__33887));
    InMux I__6553 (
            .O(N__33947),
            .I(N__33887));
    InMux I__6552 (
            .O(N__33946),
            .I(N__33887));
    InMux I__6551 (
            .O(N__33945),
            .I(N__33887));
    Span4Mux_v I__6550 (
            .O(N__33942),
            .I(N__33884));
    Span4Mux_h I__6549 (
            .O(N__33937),
            .I(N__33881));
    InMux I__6548 (
            .O(N__33936),
            .I(N__33878));
    InMux I__6547 (
            .O(N__33935),
            .I(N__33867));
    InMux I__6546 (
            .O(N__33932),
            .I(N__33867));
    InMux I__6545 (
            .O(N__33929),
            .I(N__33867));
    InMux I__6544 (
            .O(N__33928),
            .I(N__33867));
    InMux I__6543 (
            .O(N__33927),
            .I(N__33867));
    InMux I__6542 (
            .O(N__33924),
            .I(N__33858));
    InMux I__6541 (
            .O(N__33923),
            .I(N__33858));
    InMux I__6540 (
            .O(N__33922),
            .I(N__33858));
    InMux I__6539 (
            .O(N__33921),
            .I(N__33858));
    InMux I__6538 (
            .O(N__33918),
            .I(N__33841));
    InMux I__6537 (
            .O(N__33915),
            .I(N__33841));
    InMux I__6536 (
            .O(N__33912),
            .I(N__33841));
    InMux I__6535 (
            .O(N__33911),
            .I(N__33841));
    InMux I__6534 (
            .O(N__33910),
            .I(N__33841));
    InMux I__6533 (
            .O(N__33909),
            .I(N__33841));
    InMux I__6532 (
            .O(N__33908),
            .I(N__33841));
    InMux I__6531 (
            .O(N__33907),
            .I(N__33841));
    LocalMux I__6530 (
            .O(N__33904),
            .I(N__33836));
    LocalMux I__6529 (
            .O(N__33887),
            .I(N__33836));
    Span4Mux_h I__6528 (
            .O(N__33884),
            .I(N__33831));
    Span4Mux_h I__6527 (
            .O(N__33881),
            .I(N__33831));
    LocalMux I__6526 (
            .O(N__33878),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__6525 (
            .O(N__33867),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__6524 (
            .O(N__33858),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__6523 (
            .O(N__33841),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv12 I__6522 (
            .O(N__33836),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__6521 (
            .O(N__33831),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__6520 (
            .O(N__33818),
            .I(N__33815));
    InMux I__6519 (
            .O(N__33815),
            .I(N__33812));
    LocalMux I__6518 (
            .O(N__33812),
            .I(N__33809));
    Span4Mux_v I__6517 (
            .O(N__33809),
            .I(N__33806));
    Odrv4 I__6516 (
            .O(N__33806),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__6515 (
            .O(N__33803),
            .I(N__33800));
    LocalMux I__6514 (
            .O(N__33800),
            .I(N__33795));
    InMux I__6513 (
            .O(N__33799),
            .I(N__33790));
    InMux I__6512 (
            .O(N__33798),
            .I(N__33790));
    Span12Mux_h I__6511 (
            .O(N__33795),
            .I(N__33787));
    LocalMux I__6510 (
            .O(N__33790),
            .I(N__33784));
    Span12Mux_v I__6509 (
            .O(N__33787),
            .I(N__33781));
    Span12Mux_v I__6508 (
            .O(N__33784),
            .I(N__33778));
    Odrv12 I__6507 (
            .O(N__33781),
            .I(il_max_comp1_D2));
    Odrv12 I__6506 (
            .O(N__33778),
            .I(il_max_comp1_D2));
    InMux I__6505 (
            .O(N__33773),
            .I(N__33770));
    LocalMux I__6504 (
            .O(N__33770),
            .I(N__33766));
    InMux I__6503 (
            .O(N__33769),
            .I(N__33763));
    Span4Mux_h I__6502 (
            .O(N__33766),
            .I(N__33758));
    LocalMux I__6501 (
            .O(N__33763),
            .I(N__33758));
    Odrv4 I__6500 (
            .O(N__33758),
            .I(state_ns_i_a3_1));
    InMux I__6499 (
            .O(N__33755),
            .I(N__33752));
    LocalMux I__6498 (
            .O(N__33752),
            .I(N__33747));
    InMux I__6497 (
            .O(N__33751),
            .I(N__33744));
    InMux I__6496 (
            .O(N__33750),
            .I(N__33740));
    Span4Mux_v I__6495 (
            .O(N__33747),
            .I(N__33735));
    LocalMux I__6494 (
            .O(N__33744),
            .I(N__33735));
    InMux I__6493 (
            .O(N__33743),
            .I(N__33732));
    LocalMux I__6492 (
            .O(N__33740),
            .I(N__33729));
    Span4Mux_v I__6491 (
            .O(N__33735),
            .I(N__33725));
    LocalMux I__6490 (
            .O(N__33732),
            .I(N__33720));
    Span4Mux_h I__6489 (
            .O(N__33729),
            .I(N__33720));
    InMux I__6488 (
            .O(N__33728),
            .I(N__33717));
    Span4Mux_h I__6487 (
            .O(N__33725),
            .I(N__33714));
    Span4Mux_v I__6486 (
            .O(N__33720),
            .I(N__33711));
    LocalMux I__6485 (
            .O(N__33717),
            .I(measured_delay_hc_12));
    Odrv4 I__6484 (
            .O(N__33714),
            .I(measured_delay_hc_12));
    Odrv4 I__6483 (
            .O(N__33711),
            .I(measured_delay_hc_12));
    InMux I__6482 (
            .O(N__33704),
            .I(N__33699));
    InMux I__6481 (
            .O(N__33703),
            .I(N__33695));
    InMux I__6480 (
            .O(N__33702),
            .I(N__33692));
    LocalMux I__6479 (
            .O(N__33699),
            .I(N__33689));
    InMux I__6478 (
            .O(N__33698),
            .I(N__33686));
    LocalMux I__6477 (
            .O(N__33695),
            .I(N__33682));
    LocalMux I__6476 (
            .O(N__33692),
            .I(N__33679));
    Span4Mux_h I__6475 (
            .O(N__33689),
            .I(N__33674));
    LocalMux I__6474 (
            .O(N__33686),
            .I(N__33674));
    InMux I__6473 (
            .O(N__33685),
            .I(N__33671));
    Span4Mux_h I__6472 (
            .O(N__33682),
            .I(N__33668));
    Span4Mux_v I__6471 (
            .O(N__33679),
            .I(N__33665));
    Span4Mux_h I__6470 (
            .O(N__33674),
            .I(N__33662));
    LocalMux I__6469 (
            .O(N__33671),
            .I(N__33659));
    Span4Mux_v I__6468 (
            .O(N__33668),
            .I(N__33654));
    Span4Mux_h I__6467 (
            .O(N__33665),
            .I(N__33654));
    Span4Mux_v I__6466 (
            .O(N__33662),
            .I(N__33651));
    Odrv4 I__6465 (
            .O(N__33659),
            .I(measured_delay_hc_11));
    Odrv4 I__6464 (
            .O(N__33654),
            .I(measured_delay_hc_11));
    Odrv4 I__6463 (
            .O(N__33651),
            .I(measured_delay_hc_11));
    CascadeMux I__6462 (
            .O(N__33644),
            .I(N__33639));
    InMux I__6461 (
            .O(N__33643),
            .I(N__33636));
    CascadeMux I__6460 (
            .O(N__33642),
            .I(N__33632));
    InMux I__6459 (
            .O(N__33639),
            .I(N__33629));
    LocalMux I__6458 (
            .O(N__33636),
            .I(N__33626));
    InMux I__6457 (
            .O(N__33635),
            .I(N__33623));
    InMux I__6456 (
            .O(N__33632),
            .I(N__33620));
    LocalMux I__6455 (
            .O(N__33629),
            .I(N__33616));
    Span4Mux_v I__6454 (
            .O(N__33626),
            .I(N__33611));
    LocalMux I__6453 (
            .O(N__33623),
            .I(N__33611));
    LocalMux I__6452 (
            .O(N__33620),
            .I(N__33608));
    InMux I__6451 (
            .O(N__33619),
            .I(N__33605));
    Span4Mux_v I__6450 (
            .O(N__33616),
            .I(N__33598));
    Span4Mux_v I__6449 (
            .O(N__33611),
            .I(N__33598));
    Span4Mux_v I__6448 (
            .O(N__33608),
            .I(N__33598));
    LocalMux I__6447 (
            .O(N__33605),
            .I(measured_delay_hc_9));
    Odrv4 I__6446 (
            .O(N__33598),
            .I(measured_delay_hc_9));
    CascadeMux I__6445 (
            .O(N__33593),
            .I(N__33589));
    CascadeMux I__6444 (
            .O(N__33592),
            .I(N__33586));
    InMux I__6443 (
            .O(N__33589),
            .I(N__33582));
    InMux I__6442 (
            .O(N__33586),
            .I(N__33578));
    InMux I__6441 (
            .O(N__33585),
            .I(N__33575));
    LocalMux I__6440 (
            .O(N__33582),
            .I(N__33571));
    InMux I__6439 (
            .O(N__33581),
            .I(N__33568));
    LocalMux I__6438 (
            .O(N__33578),
            .I(N__33565));
    LocalMux I__6437 (
            .O(N__33575),
            .I(N__33562));
    InMux I__6436 (
            .O(N__33574),
            .I(N__33559));
    Span4Mux_v I__6435 (
            .O(N__33571),
            .I(N__33556));
    LocalMux I__6434 (
            .O(N__33568),
            .I(N__33553));
    Span4Mux_v I__6433 (
            .O(N__33565),
            .I(N__33548));
    Span4Mux_v I__6432 (
            .O(N__33562),
            .I(N__33548));
    LocalMux I__6431 (
            .O(N__33559),
            .I(N__33545));
    Span4Mux_h I__6430 (
            .O(N__33556),
            .I(N__33540));
    Span4Mux_v I__6429 (
            .O(N__33553),
            .I(N__33540));
    Odrv4 I__6428 (
            .O(N__33548),
            .I(measured_delay_hc_10));
    Odrv12 I__6427 (
            .O(N__33545),
            .I(measured_delay_hc_10));
    Odrv4 I__6426 (
            .O(N__33540),
            .I(measured_delay_hc_10));
    InMux I__6425 (
            .O(N__33533),
            .I(N__33530));
    LocalMux I__6424 (
            .O(N__33530),
            .I(N__33527));
    Odrv4 I__6423 (
            .O(N__33527),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ));
    InMux I__6422 (
            .O(N__33524),
            .I(N__33504));
    CascadeMux I__6421 (
            .O(N__33523),
            .I(N__33501));
    CascadeMux I__6420 (
            .O(N__33522),
            .I(N__33496));
    InMux I__6419 (
            .O(N__33521),
            .I(N__33491));
    InMux I__6418 (
            .O(N__33520),
            .I(N__33491));
    InMux I__6417 (
            .O(N__33519),
            .I(N__33482));
    InMux I__6416 (
            .O(N__33518),
            .I(N__33482));
    InMux I__6415 (
            .O(N__33517),
            .I(N__33482));
    InMux I__6414 (
            .O(N__33516),
            .I(N__33482));
    InMux I__6413 (
            .O(N__33515),
            .I(N__33479));
    InMux I__6412 (
            .O(N__33514),
            .I(N__33470));
    InMux I__6411 (
            .O(N__33513),
            .I(N__33465));
    InMux I__6410 (
            .O(N__33512),
            .I(N__33465));
    InMux I__6409 (
            .O(N__33511),
            .I(N__33460));
    InMux I__6408 (
            .O(N__33510),
            .I(N__33460));
    InMux I__6407 (
            .O(N__33509),
            .I(N__33453));
    InMux I__6406 (
            .O(N__33508),
            .I(N__33453));
    InMux I__6405 (
            .O(N__33507),
            .I(N__33453));
    LocalMux I__6404 (
            .O(N__33504),
            .I(N__33448));
    InMux I__6403 (
            .O(N__33501),
            .I(N__33443));
    InMux I__6402 (
            .O(N__33500),
            .I(N__33443));
    InMux I__6401 (
            .O(N__33499),
            .I(N__33438));
    InMux I__6400 (
            .O(N__33496),
            .I(N__33438));
    LocalMux I__6399 (
            .O(N__33491),
            .I(N__33432));
    LocalMux I__6398 (
            .O(N__33482),
            .I(N__33432));
    LocalMux I__6397 (
            .O(N__33479),
            .I(N__33429));
    InMux I__6396 (
            .O(N__33478),
            .I(N__33418));
    InMux I__6395 (
            .O(N__33477),
            .I(N__33418));
    InMux I__6394 (
            .O(N__33476),
            .I(N__33418));
    InMux I__6393 (
            .O(N__33475),
            .I(N__33418));
    InMux I__6392 (
            .O(N__33474),
            .I(N__33418));
    InMux I__6391 (
            .O(N__33473),
            .I(N__33415));
    LocalMux I__6390 (
            .O(N__33470),
            .I(N__33411));
    LocalMux I__6389 (
            .O(N__33465),
            .I(N__33408));
    LocalMux I__6388 (
            .O(N__33460),
            .I(N__33405));
    LocalMux I__6387 (
            .O(N__33453),
            .I(N__33402));
    InMux I__6386 (
            .O(N__33452),
            .I(N__33397));
    InMux I__6385 (
            .O(N__33451),
            .I(N__33397));
    Span4Mux_v I__6384 (
            .O(N__33448),
            .I(N__33392));
    LocalMux I__6383 (
            .O(N__33443),
            .I(N__33392));
    LocalMux I__6382 (
            .O(N__33438),
            .I(N__33389));
    InMux I__6381 (
            .O(N__33437),
            .I(N__33386));
    Span4Mux_v I__6380 (
            .O(N__33432),
            .I(N__33379));
    Span4Mux_h I__6379 (
            .O(N__33429),
            .I(N__33379));
    LocalMux I__6378 (
            .O(N__33418),
            .I(N__33379));
    LocalMux I__6377 (
            .O(N__33415),
            .I(N__33373));
    InMux I__6376 (
            .O(N__33414),
            .I(N__33370));
    Span4Mux_v I__6375 (
            .O(N__33411),
            .I(N__33359));
    Span4Mux_v I__6374 (
            .O(N__33408),
            .I(N__33359));
    Span4Mux_v I__6373 (
            .O(N__33405),
            .I(N__33359));
    Span4Mux_v I__6372 (
            .O(N__33402),
            .I(N__33359));
    LocalMux I__6371 (
            .O(N__33397),
            .I(N__33359));
    Span4Mux_h I__6370 (
            .O(N__33392),
            .I(N__33354));
    Span4Mux_h I__6369 (
            .O(N__33389),
            .I(N__33354));
    LocalMux I__6368 (
            .O(N__33386),
            .I(N__33349));
    Span4Mux_h I__6367 (
            .O(N__33379),
            .I(N__33349));
    InMux I__6366 (
            .O(N__33378),
            .I(N__33344));
    InMux I__6365 (
            .O(N__33377),
            .I(N__33344));
    InMux I__6364 (
            .O(N__33376),
            .I(N__33341));
    Odrv4 I__6363 (
            .O(N__33373),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__6362 (
            .O(N__33370),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__6361 (
            .O(N__33359),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__6360 (
            .O(N__33354),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__6359 (
            .O(N__33349),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__6358 (
            .O(N__33344),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__6357 (
            .O(N__33341),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    CascadeMux I__6356 (
            .O(N__33326),
            .I(N__33309));
    InMux I__6355 (
            .O(N__33325),
            .I(N__33302));
    InMux I__6354 (
            .O(N__33324),
            .I(N__33302));
    InMux I__6353 (
            .O(N__33323),
            .I(N__33297));
    InMux I__6352 (
            .O(N__33322),
            .I(N__33297));
    InMux I__6351 (
            .O(N__33321),
            .I(N__33294));
    InMux I__6350 (
            .O(N__33320),
            .I(N__33290));
    InMux I__6349 (
            .O(N__33319),
            .I(N__33286));
    InMux I__6348 (
            .O(N__33318),
            .I(N__33283));
    InMux I__6347 (
            .O(N__33317),
            .I(N__33280));
    InMux I__6346 (
            .O(N__33316),
            .I(N__33277));
    InMux I__6345 (
            .O(N__33315),
            .I(N__33274));
    InMux I__6344 (
            .O(N__33314),
            .I(N__33268));
    InMux I__6343 (
            .O(N__33313),
            .I(N__33263));
    InMux I__6342 (
            .O(N__33312),
            .I(N__33263));
    InMux I__6341 (
            .O(N__33309),
            .I(N__33252));
    InMux I__6340 (
            .O(N__33308),
            .I(N__33252));
    InMux I__6339 (
            .O(N__33307),
            .I(N__33252));
    LocalMux I__6338 (
            .O(N__33302),
            .I(N__33245));
    LocalMux I__6337 (
            .O(N__33297),
            .I(N__33245));
    LocalMux I__6336 (
            .O(N__33294),
            .I(N__33245));
    InMux I__6335 (
            .O(N__33293),
            .I(N__33242));
    LocalMux I__6334 (
            .O(N__33290),
            .I(N__33239));
    InMux I__6333 (
            .O(N__33289),
            .I(N__33236));
    LocalMux I__6332 (
            .O(N__33286),
            .I(N__33231));
    LocalMux I__6331 (
            .O(N__33283),
            .I(N__33231));
    LocalMux I__6330 (
            .O(N__33280),
            .I(N__33224));
    LocalMux I__6329 (
            .O(N__33277),
            .I(N__33224));
    LocalMux I__6328 (
            .O(N__33274),
            .I(N__33224));
    InMux I__6327 (
            .O(N__33273),
            .I(N__33217));
    InMux I__6326 (
            .O(N__33272),
            .I(N__33217));
    InMux I__6325 (
            .O(N__33271),
            .I(N__33217));
    LocalMux I__6324 (
            .O(N__33268),
            .I(N__33212));
    LocalMux I__6323 (
            .O(N__33263),
            .I(N__33212));
    InMux I__6322 (
            .O(N__33262),
            .I(N__33207));
    InMux I__6321 (
            .O(N__33261),
            .I(N__33207));
    InMux I__6320 (
            .O(N__33260),
            .I(N__33197));
    InMux I__6319 (
            .O(N__33259),
            .I(N__33197));
    LocalMux I__6318 (
            .O(N__33252),
            .I(N__33188));
    Span4Mux_v I__6317 (
            .O(N__33245),
            .I(N__33188));
    LocalMux I__6316 (
            .O(N__33242),
            .I(N__33188));
    Span4Mux_v I__6315 (
            .O(N__33239),
            .I(N__33188));
    LocalMux I__6314 (
            .O(N__33236),
            .I(N__33185));
    Span4Mux_h I__6313 (
            .O(N__33231),
            .I(N__33180));
    Span4Mux_v I__6312 (
            .O(N__33224),
            .I(N__33180));
    LocalMux I__6311 (
            .O(N__33217),
            .I(N__33177));
    Span4Mux_h I__6310 (
            .O(N__33212),
            .I(N__33172));
    LocalMux I__6309 (
            .O(N__33207),
            .I(N__33172));
    InMux I__6308 (
            .O(N__33206),
            .I(N__33163));
    InMux I__6307 (
            .O(N__33205),
            .I(N__33163));
    InMux I__6306 (
            .O(N__33204),
            .I(N__33163));
    InMux I__6305 (
            .O(N__33203),
            .I(N__33163));
    InMux I__6304 (
            .O(N__33202),
            .I(N__33160));
    LocalMux I__6303 (
            .O(N__33197),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6302 (
            .O(N__33188),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6301 (
            .O(N__33185),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6300 (
            .O(N__33180),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6299 (
            .O(N__33177),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6298 (
            .O(N__33172),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__6297 (
            .O(N__33163),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__6296 (
            .O(N__33160),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    InMux I__6295 (
            .O(N__33143),
            .I(N__33133));
    InMux I__6294 (
            .O(N__33142),
            .I(N__33124));
    InMux I__6293 (
            .O(N__33141),
            .I(N__33119));
    InMux I__6292 (
            .O(N__33140),
            .I(N__33114));
    InMux I__6291 (
            .O(N__33139),
            .I(N__33114));
    InMux I__6290 (
            .O(N__33138),
            .I(N__33107));
    InMux I__6289 (
            .O(N__33137),
            .I(N__33107));
    InMux I__6288 (
            .O(N__33136),
            .I(N__33107));
    LocalMux I__6287 (
            .O(N__33133),
            .I(N__33104));
    InMux I__6286 (
            .O(N__33132),
            .I(N__33099));
    InMux I__6285 (
            .O(N__33131),
            .I(N__33099));
    InMux I__6284 (
            .O(N__33130),
            .I(N__33094));
    InMux I__6283 (
            .O(N__33129),
            .I(N__33094));
    InMux I__6282 (
            .O(N__33128),
            .I(N__33091));
    InMux I__6281 (
            .O(N__33127),
            .I(N__33086));
    LocalMux I__6280 (
            .O(N__33124),
            .I(N__33083));
    InMux I__6279 (
            .O(N__33123),
            .I(N__33078));
    InMux I__6278 (
            .O(N__33122),
            .I(N__33078));
    LocalMux I__6277 (
            .O(N__33119),
            .I(N__33072));
    LocalMux I__6276 (
            .O(N__33114),
            .I(N__33069));
    LocalMux I__6275 (
            .O(N__33107),
            .I(N__33060));
    Span4Mux_h I__6274 (
            .O(N__33104),
            .I(N__33060));
    LocalMux I__6273 (
            .O(N__33099),
            .I(N__33060));
    LocalMux I__6272 (
            .O(N__33094),
            .I(N__33060));
    LocalMux I__6271 (
            .O(N__33091),
            .I(N__33055));
    InMux I__6270 (
            .O(N__33090),
            .I(N__33050));
    InMux I__6269 (
            .O(N__33089),
            .I(N__33050));
    LocalMux I__6268 (
            .O(N__33086),
            .I(N__33038));
    Span4Mux_h I__6267 (
            .O(N__33083),
            .I(N__33033));
    LocalMux I__6266 (
            .O(N__33078),
            .I(N__33033));
    InMux I__6265 (
            .O(N__33077),
            .I(N__33030));
    InMux I__6264 (
            .O(N__33076),
            .I(N__33025));
    InMux I__6263 (
            .O(N__33075),
            .I(N__33025));
    Span4Mux_h I__6262 (
            .O(N__33072),
            .I(N__33018));
    Span4Mux_v I__6261 (
            .O(N__33069),
            .I(N__33018));
    Span4Mux_v I__6260 (
            .O(N__33060),
            .I(N__33018));
    InMux I__6259 (
            .O(N__33059),
            .I(N__33013));
    InMux I__6258 (
            .O(N__33058),
            .I(N__33013));
    Span4Mux_h I__6257 (
            .O(N__33055),
            .I(N__33008));
    LocalMux I__6256 (
            .O(N__33050),
            .I(N__33008));
    InMux I__6255 (
            .O(N__33049),
            .I(N__32999));
    InMux I__6254 (
            .O(N__33048),
            .I(N__32999));
    InMux I__6253 (
            .O(N__33047),
            .I(N__32999));
    InMux I__6252 (
            .O(N__33046),
            .I(N__32999));
    InMux I__6251 (
            .O(N__33045),
            .I(N__32988));
    InMux I__6250 (
            .O(N__33044),
            .I(N__32988));
    InMux I__6249 (
            .O(N__33043),
            .I(N__32988));
    InMux I__6248 (
            .O(N__33042),
            .I(N__32988));
    InMux I__6247 (
            .O(N__33041),
            .I(N__32988));
    Odrv4 I__6246 (
            .O(N__33038),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    Odrv4 I__6245 (
            .O(N__33033),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    LocalMux I__6244 (
            .O(N__33030),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    LocalMux I__6243 (
            .O(N__33025),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    Odrv4 I__6242 (
            .O(N__33018),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    LocalMux I__6241 (
            .O(N__33013),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    Odrv4 I__6240 (
            .O(N__33008),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    LocalMux I__6239 (
            .O(N__32999),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    LocalMux I__6238 (
            .O(N__32988),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    InMux I__6237 (
            .O(N__32969),
            .I(N__32964));
    InMux I__6236 (
            .O(N__32968),
            .I(N__32961));
    CascadeMux I__6235 (
            .O(N__32967),
            .I(N__32958));
    LocalMux I__6234 (
            .O(N__32964),
            .I(N__32955));
    LocalMux I__6233 (
            .O(N__32961),
            .I(N__32952));
    InMux I__6232 (
            .O(N__32958),
            .I(N__32949));
    Sp12to4 I__6231 (
            .O(N__32955),
            .I(N__32946));
    Span4Mux_h I__6230 (
            .O(N__32952),
            .I(N__32943));
    LocalMux I__6229 (
            .O(N__32949),
            .I(measured_delay_hc_22));
    Odrv12 I__6228 (
            .O(N__32946),
            .I(measured_delay_hc_22));
    Odrv4 I__6227 (
            .O(N__32943),
            .I(measured_delay_hc_22));
    CascadeMux I__6226 (
            .O(N__32936),
            .I(N__32931));
    InMux I__6225 (
            .O(N__32935),
            .I(N__32928));
    InMux I__6224 (
            .O(N__32934),
            .I(N__32924));
    InMux I__6223 (
            .O(N__32931),
            .I(N__32921));
    LocalMux I__6222 (
            .O(N__32928),
            .I(N__32917));
    InMux I__6221 (
            .O(N__32927),
            .I(N__32914));
    LocalMux I__6220 (
            .O(N__32924),
            .I(N__32909));
    LocalMux I__6219 (
            .O(N__32921),
            .I(N__32909));
    CascadeMux I__6218 (
            .O(N__32920),
            .I(N__32906));
    Span4Mux_v I__6217 (
            .O(N__32917),
            .I(N__32899));
    LocalMux I__6216 (
            .O(N__32914),
            .I(N__32899));
    Span4Mux_h I__6215 (
            .O(N__32909),
            .I(N__32899));
    InMux I__6214 (
            .O(N__32906),
            .I(N__32896));
    Span4Mux_h I__6213 (
            .O(N__32899),
            .I(N__32893));
    LocalMux I__6212 (
            .O(N__32896),
            .I(measured_delay_hc_16));
    Odrv4 I__6211 (
            .O(N__32893),
            .I(measured_delay_hc_16));
    CascadeMux I__6210 (
            .O(N__32888),
            .I(N__32885));
    InMux I__6209 (
            .O(N__32885),
            .I(N__32882));
    LocalMux I__6208 (
            .O(N__32882),
            .I(N__32879));
    Odrv4 I__6207 (
            .O(N__32879),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__6206 (
            .O(N__32876),
            .I(N__32872));
    InMux I__6205 (
            .O(N__32875),
            .I(N__32867));
    LocalMux I__6204 (
            .O(N__32872),
            .I(N__32863));
    InMux I__6203 (
            .O(N__32871),
            .I(N__32858));
    InMux I__6202 (
            .O(N__32870),
            .I(N__32858));
    LocalMux I__6201 (
            .O(N__32867),
            .I(N__32855));
    InMux I__6200 (
            .O(N__32866),
            .I(N__32852));
    Span4Mux_h I__6199 (
            .O(N__32863),
            .I(N__32847));
    LocalMux I__6198 (
            .O(N__32858),
            .I(N__32847));
    Span12Mux_s11_h I__6197 (
            .O(N__32855),
            .I(N__32844));
    LocalMux I__6196 (
            .O(N__32852),
            .I(N__32841));
    Span4Mux_v I__6195 (
            .O(N__32847),
            .I(N__32838));
    Odrv12 I__6194 (
            .O(N__32844),
            .I(measured_delay_hc_1));
    Odrv4 I__6193 (
            .O(N__32841),
            .I(measured_delay_hc_1));
    Odrv4 I__6192 (
            .O(N__32838),
            .I(measured_delay_hc_1));
    CascadeMux I__6191 (
            .O(N__32831),
            .I(N__32828));
    InMux I__6190 (
            .O(N__32828),
            .I(N__32825));
    LocalMux I__6189 (
            .O(N__32825),
            .I(N__32822));
    Odrv12 I__6188 (
            .O(N__32822),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    InMux I__6187 (
            .O(N__32819),
            .I(N__32811));
    InMux I__6186 (
            .O(N__32818),
            .I(N__32811));
    InMux I__6185 (
            .O(N__32817),
            .I(N__32806));
    InMux I__6184 (
            .O(N__32816),
            .I(N__32806));
    LocalMux I__6183 (
            .O(N__32811),
            .I(N__32803));
    LocalMux I__6182 (
            .O(N__32806),
            .I(N__32800));
    Odrv4 I__6181 (
            .O(N__32803),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    Odrv12 I__6180 (
            .O(N__32800),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    InMux I__6179 (
            .O(N__32795),
            .I(N__32791));
    InMux I__6178 (
            .O(N__32794),
            .I(N__32785));
    LocalMux I__6177 (
            .O(N__32791),
            .I(N__32782));
    InMux I__6176 (
            .O(N__32790),
            .I(N__32779));
    CascadeMux I__6175 (
            .O(N__32789),
            .I(N__32776));
    CascadeMux I__6174 (
            .O(N__32788),
            .I(N__32773));
    LocalMux I__6173 (
            .O(N__32785),
            .I(N__32770));
    Span4Mux_h I__6172 (
            .O(N__32782),
            .I(N__32767));
    LocalMux I__6171 (
            .O(N__32779),
            .I(N__32764));
    InMux I__6170 (
            .O(N__32776),
            .I(N__32759));
    InMux I__6169 (
            .O(N__32773),
            .I(N__32759));
    Span4Mux_v I__6168 (
            .O(N__32770),
            .I(N__32756));
    Span4Mux_v I__6167 (
            .O(N__32767),
            .I(N__32749));
    Span4Mux_h I__6166 (
            .O(N__32764),
            .I(N__32749));
    LocalMux I__6165 (
            .O(N__32759),
            .I(N__32749));
    Odrv4 I__6164 (
            .O(N__32756),
            .I(measured_delay_hc_3));
    Odrv4 I__6163 (
            .O(N__32749),
            .I(measured_delay_hc_3));
    CascadeMux I__6162 (
            .O(N__32744),
            .I(N__32741));
    InMux I__6161 (
            .O(N__32741),
            .I(N__32738));
    LocalMux I__6160 (
            .O(N__32738),
            .I(N__32735));
    Odrv12 I__6159 (
            .O(N__32735),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__6158 (
            .O(N__32732),
            .I(N__32729));
    LocalMux I__6157 (
            .O(N__32729),
            .I(N__32726));
    Span4Mux_v I__6156 (
            .O(N__32726),
            .I(N__32720));
    InMux I__6155 (
            .O(N__32725),
            .I(N__32717));
    InMux I__6154 (
            .O(N__32724),
            .I(N__32713));
    InMux I__6153 (
            .O(N__32723),
            .I(N__32710));
    Sp12to4 I__6152 (
            .O(N__32720),
            .I(N__32705));
    LocalMux I__6151 (
            .O(N__32717),
            .I(N__32705));
    InMux I__6150 (
            .O(N__32716),
            .I(N__32702));
    LocalMux I__6149 (
            .O(N__32713),
            .I(measured_delay_hc_7));
    LocalMux I__6148 (
            .O(N__32710),
            .I(measured_delay_hc_7));
    Odrv12 I__6147 (
            .O(N__32705),
            .I(measured_delay_hc_7));
    LocalMux I__6146 (
            .O(N__32702),
            .I(measured_delay_hc_7));
    CascadeMux I__6145 (
            .O(N__32693),
            .I(N__32690));
    InMux I__6144 (
            .O(N__32690),
            .I(N__32687));
    LocalMux I__6143 (
            .O(N__32687),
            .I(N__32684));
    Span4Mux_v I__6142 (
            .O(N__32684),
            .I(N__32681));
    Odrv4 I__6141 (
            .O(N__32681),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__6140 (
            .O(N__32678),
            .I(N__32675));
    LocalMux I__6139 (
            .O(N__32675),
            .I(N__32671));
    InMux I__6138 (
            .O(N__32674),
            .I(N__32667));
    Span4Mux_h I__6137 (
            .O(N__32671),
            .I(N__32663));
    InMux I__6136 (
            .O(N__32670),
            .I(N__32660));
    LocalMux I__6135 (
            .O(N__32667),
            .I(N__32656));
    InMux I__6134 (
            .O(N__32666),
            .I(N__32653));
    Span4Mux_v I__6133 (
            .O(N__32663),
            .I(N__32650));
    LocalMux I__6132 (
            .O(N__32660),
            .I(N__32647));
    InMux I__6131 (
            .O(N__32659),
            .I(N__32644));
    Span4Mux_h I__6130 (
            .O(N__32656),
            .I(N__32639));
    LocalMux I__6129 (
            .O(N__32653),
            .I(N__32639));
    Span4Mux_h I__6128 (
            .O(N__32650),
            .I(N__32636));
    Span4Mux_v I__6127 (
            .O(N__32647),
            .I(N__32631));
    LocalMux I__6126 (
            .O(N__32644),
            .I(N__32631));
    Span4Mux_h I__6125 (
            .O(N__32639),
            .I(N__32628));
    Odrv4 I__6124 (
            .O(N__32636),
            .I(measured_delay_hc_8));
    Odrv4 I__6123 (
            .O(N__32631),
            .I(measured_delay_hc_8));
    Odrv4 I__6122 (
            .O(N__32628),
            .I(measured_delay_hc_8));
    CascadeMux I__6121 (
            .O(N__32621),
            .I(N__32618));
    InMux I__6120 (
            .O(N__32618),
            .I(N__32615));
    LocalMux I__6119 (
            .O(N__32615),
            .I(N__32612));
    Odrv12 I__6118 (
            .O(N__32612),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__6117 (
            .O(N__32609),
            .I(N__32606));
    InMux I__6116 (
            .O(N__32606),
            .I(N__32603));
    LocalMux I__6115 (
            .O(N__32603),
            .I(N__32600));
    Span4Mux_h I__6114 (
            .O(N__32600),
            .I(N__32597));
    Odrv4 I__6113 (
            .O(N__32597),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__6112 (
            .O(N__32594),
            .I(N__32591));
    InMux I__6111 (
            .O(N__32591),
            .I(N__32588));
    LocalMux I__6110 (
            .O(N__32588),
            .I(N__32585));
    Span4Mux_h I__6109 (
            .O(N__32585),
            .I(N__32582));
    Odrv4 I__6108 (
            .O(N__32582),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__6107 (
            .O(N__32579),
            .I(N__32576));
    LocalMux I__6106 (
            .O(N__32576),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13 ));
    CascadeMux I__6105 (
            .O(N__32573),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ));
    InMux I__6104 (
            .O(N__32570),
            .I(N__32566));
    InMux I__6103 (
            .O(N__32569),
            .I(N__32562));
    LocalMux I__6102 (
            .O(N__32566),
            .I(N__32559));
    InMux I__6101 (
            .O(N__32565),
            .I(N__32555));
    LocalMux I__6100 (
            .O(N__32562),
            .I(N__32552));
    Span4Mux_v I__6099 (
            .O(N__32559),
            .I(N__32549));
    InMux I__6098 (
            .O(N__32558),
            .I(N__32546));
    LocalMux I__6097 (
            .O(N__32555),
            .I(measured_delay_hc_0));
    Odrv12 I__6096 (
            .O(N__32552),
            .I(measured_delay_hc_0));
    Odrv4 I__6095 (
            .O(N__32549),
            .I(measured_delay_hc_0));
    LocalMux I__6094 (
            .O(N__32546),
            .I(measured_delay_hc_0));
    InMux I__6093 (
            .O(N__32537),
            .I(N__32534));
    LocalMux I__6092 (
            .O(N__32534),
            .I(N__32531));
    Odrv12 I__6091 (
            .O(N__32531),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ));
    InMux I__6090 (
            .O(N__32528),
            .I(N__32525));
    LocalMux I__6089 (
            .O(N__32525),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__6088 (
            .O(N__32522),
            .I(N__32518));
    InMux I__6087 (
            .O(N__32521),
            .I(N__32515));
    LocalMux I__6086 (
            .O(N__32518),
            .I(N__32512));
    LocalMux I__6085 (
            .O(N__32515),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__6084 (
            .O(N__32512),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__6083 (
            .O(N__32507),
            .I(N__32504));
    LocalMux I__6082 (
            .O(N__32504),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__6081 (
            .O(N__32501),
            .I(N__32497));
    InMux I__6080 (
            .O(N__32500),
            .I(N__32494));
    LocalMux I__6079 (
            .O(N__32497),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__6078 (
            .O(N__32494),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__6077 (
            .O(N__32489),
            .I(N__32486));
    LocalMux I__6076 (
            .O(N__32486),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__6075 (
            .O(N__32483),
            .I(N__32479));
    InMux I__6074 (
            .O(N__32482),
            .I(N__32476));
    LocalMux I__6073 (
            .O(N__32479),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__6072 (
            .O(N__32476),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__6071 (
            .O(N__32471),
            .I(N__32468));
    LocalMux I__6070 (
            .O(N__32468),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__6069 (
            .O(N__32465),
            .I(N__32461));
    InMux I__6068 (
            .O(N__32464),
            .I(N__32458));
    LocalMux I__6067 (
            .O(N__32461),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__6066 (
            .O(N__32458),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__6065 (
            .O(N__32453),
            .I(N__32450));
    LocalMux I__6064 (
            .O(N__32450),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__6063 (
            .O(N__32447),
            .I(N__32443));
    InMux I__6062 (
            .O(N__32446),
            .I(N__32440));
    LocalMux I__6061 (
            .O(N__32443),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__6060 (
            .O(N__32440),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__6059 (
            .O(N__32435),
            .I(N__32432));
    LocalMux I__6058 (
            .O(N__32432),
            .I(N__32427));
    InMux I__6057 (
            .O(N__32431),
            .I(N__32422));
    InMux I__6056 (
            .O(N__32430),
            .I(N__32419));
    Span4Mux_v I__6055 (
            .O(N__32427),
            .I(N__32416));
    InMux I__6054 (
            .O(N__32426),
            .I(N__32413));
    InMux I__6053 (
            .O(N__32425),
            .I(N__32410));
    LocalMux I__6052 (
            .O(N__32422),
            .I(N__32407));
    LocalMux I__6051 (
            .O(N__32419),
            .I(N__32404));
    Span4Mux_v I__6050 (
            .O(N__32416),
            .I(N__32401));
    LocalMux I__6049 (
            .O(N__32413),
            .I(N__32398));
    LocalMux I__6048 (
            .O(N__32410),
            .I(N__32395));
    Span4Mux_h I__6047 (
            .O(N__32407),
            .I(N__32390));
    Span4Mux_h I__6046 (
            .O(N__32404),
            .I(N__32390));
    Odrv4 I__6045 (
            .O(N__32401),
            .I(measured_delay_hc_4));
    Odrv12 I__6044 (
            .O(N__32398),
            .I(measured_delay_hc_4));
    Odrv4 I__6043 (
            .O(N__32395),
            .I(measured_delay_hc_4));
    Odrv4 I__6042 (
            .O(N__32390),
            .I(measured_delay_hc_4));
    CascadeMux I__6041 (
            .O(N__32381),
            .I(N__32378));
    InMux I__6040 (
            .O(N__32378),
            .I(N__32375));
    LocalMux I__6039 (
            .O(N__32375),
            .I(N__32372));
    Odrv12 I__6038 (
            .O(N__32372),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    InMux I__6037 (
            .O(N__32369),
            .I(N__32366));
    LocalMux I__6036 (
            .O(N__32366),
            .I(N__32361));
    InMux I__6035 (
            .O(N__32365),
            .I(N__32358));
    InMux I__6034 (
            .O(N__32364),
            .I(N__32353));
    Span4Mux_v I__6033 (
            .O(N__32361),
            .I(N__32350));
    LocalMux I__6032 (
            .O(N__32358),
            .I(N__32347));
    InMux I__6031 (
            .O(N__32357),
            .I(N__32344));
    InMux I__6030 (
            .O(N__32356),
            .I(N__32341));
    LocalMux I__6029 (
            .O(N__32353),
            .I(N__32338));
    Odrv4 I__6028 (
            .O(N__32350),
            .I(measured_delay_hc_5));
    Odrv4 I__6027 (
            .O(N__32347),
            .I(measured_delay_hc_5));
    LocalMux I__6026 (
            .O(N__32344),
            .I(measured_delay_hc_5));
    LocalMux I__6025 (
            .O(N__32341),
            .I(measured_delay_hc_5));
    Odrv4 I__6024 (
            .O(N__32338),
            .I(measured_delay_hc_5));
    CascadeMux I__6023 (
            .O(N__32327),
            .I(N__32324));
    InMux I__6022 (
            .O(N__32324),
            .I(N__32321));
    LocalMux I__6021 (
            .O(N__32321),
            .I(N__32318));
    Span4Mux_h I__6020 (
            .O(N__32318),
            .I(N__32315));
    Odrv4 I__6019 (
            .O(N__32315),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__6018 (
            .O(N__32312),
            .I(N__32309));
    InMux I__6017 (
            .O(N__32309),
            .I(N__32306));
    LocalMux I__6016 (
            .O(N__32306),
            .I(N__32303));
    Span4Mux_h I__6015 (
            .O(N__32303),
            .I(N__32300));
    Odrv4 I__6014 (
            .O(N__32300),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__6013 (
            .O(N__32297),
            .I(N__32294));
    InMux I__6012 (
            .O(N__32294),
            .I(N__32291));
    LocalMux I__6011 (
            .O(N__32291),
            .I(N__32288));
    Span4Mux_h I__6010 (
            .O(N__32288),
            .I(N__32285));
    Odrv4 I__6009 (
            .O(N__32285),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__6008 (
            .O(N__32282),
            .I(N__32279));
    LocalMux I__6007 (
            .O(N__32279),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ));
    InMux I__6006 (
            .O(N__32276),
            .I(N__32273));
    LocalMux I__6005 (
            .O(N__32273),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ));
    InMux I__6004 (
            .O(N__32270),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__6003 (
            .O(N__32267),
            .I(N__32264));
    LocalMux I__6002 (
            .O(N__32264),
            .I(N__32261));
    Span4Mux_h I__6001 (
            .O(N__32261),
            .I(N__32258));
    Odrv4 I__6000 (
            .O(N__32258),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__5999 (
            .O(N__32255),
            .I(N__32252));
    LocalMux I__5998 (
            .O(N__32252),
            .I(N__32249));
    Span4Mux_v I__5997 (
            .O(N__32249),
            .I(N__32246));
    Odrv4 I__5996 (
            .O(N__32246),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__5995 (
            .O(N__32243),
            .I(N__32240));
    LocalMux I__5994 (
            .O(N__32240),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__5993 (
            .O(N__32237),
            .I(N__32233));
    InMux I__5992 (
            .O(N__32236),
            .I(N__32230));
    LocalMux I__5991 (
            .O(N__32233),
            .I(N__32227));
    LocalMux I__5990 (
            .O(N__32230),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__5989 (
            .O(N__32227),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__5988 (
            .O(N__32222),
            .I(N__32219));
    LocalMux I__5987 (
            .O(N__32219),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__5986 (
            .O(N__32216),
            .I(N__32212));
    InMux I__5985 (
            .O(N__32215),
            .I(N__32209));
    LocalMux I__5984 (
            .O(N__32212),
            .I(N__32206));
    LocalMux I__5983 (
            .O(N__32209),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__5982 (
            .O(N__32206),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__5981 (
            .O(N__32201),
            .I(N__32198));
    LocalMux I__5980 (
            .O(N__32198),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__5979 (
            .O(N__32195),
            .I(N__32191));
    InMux I__5978 (
            .O(N__32194),
            .I(N__32188));
    LocalMux I__5977 (
            .O(N__32191),
            .I(N__32185));
    LocalMux I__5976 (
            .O(N__32188),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__5975 (
            .O(N__32185),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__5974 (
            .O(N__32180),
            .I(N__32177));
    LocalMux I__5973 (
            .O(N__32177),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__5972 (
            .O(N__32174),
            .I(N__32171));
    LocalMux I__5971 (
            .O(N__32171),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__5970 (
            .O(N__32168),
            .I(N__32165));
    LocalMux I__5969 (
            .O(N__32165),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__5968 (
            .O(N__32162),
            .I(N__32159));
    LocalMux I__5967 (
            .O(N__32159),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__5966 (
            .O(N__32156),
            .I(N__32153));
    InMux I__5965 (
            .O(N__32153),
            .I(N__32150));
    LocalMux I__5964 (
            .O(N__32150),
            .I(N__32147));
    Span4Mux_h I__5963 (
            .O(N__32147),
            .I(N__32144));
    Odrv4 I__5962 (
            .O(N__32144),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__5961 (
            .O(N__32141),
            .I(N__32138));
    LocalMux I__5960 (
            .O(N__32138),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__5959 (
            .O(N__32135),
            .I(N__32132));
    LocalMux I__5958 (
            .O(N__32132),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__5957 (
            .O(N__32129),
            .I(N__32126));
    LocalMux I__5956 (
            .O(N__32126),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__5955 (
            .O(N__32123),
            .I(N__32120));
    InMux I__5954 (
            .O(N__32120),
            .I(N__32117));
    LocalMux I__5953 (
            .O(N__32117),
            .I(N__32114));
    Odrv4 I__5952 (
            .O(N__32114),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__5951 (
            .O(N__32111),
            .I(N__32108));
    LocalMux I__5950 (
            .O(N__32108),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ));
    InMux I__5949 (
            .O(N__32105),
            .I(N__32102));
    LocalMux I__5948 (
            .O(N__32102),
            .I(N__32098));
    InMux I__5947 (
            .O(N__32101),
            .I(N__32095));
    Odrv4 I__5946 (
            .O(N__32098),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__5945 (
            .O(N__32095),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__5944 (
            .O(N__32090),
            .I(N__32087));
    LocalMux I__5943 (
            .O(N__32087),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__5942 (
            .O(N__32084),
            .I(N__32081));
    InMux I__5941 (
            .O(N__32081),
            .I(N__32077));
    InMux I__5940 (
            .O(N__32080),
            .I(N__32074));
    LocalMux I__5939 (
            .O(N__32077),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__5938 (
            .O(N__32074),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__5937 (
            .O(N__32069),
            .I(N__32066));
    LocalMux I__5936 (
            .O(N__32066),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__5935 (
            .O(N__32063),
            .I(N__32059));
    InMux I__5934 (
            .O(N__32062),
            .I(N__32056));
    LocalMux I__5933 (
            .O(N__32059),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__5932 (
            .O(N__32056),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__5931 (
            .O(N__32051),
            .I(N__32048));
    LocalMux I__5930 (
            .O(N__32048),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__5929 (
            .O(N__32045),
            .I(N__32041));
    InMux I__5928 (
            .O(N__32044),
            .I(N__32038));
    LocalMux I__5927 (
            .O(N__32041),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__5926 (
            .O(N__32038),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__5925 (
            .O(N__32033),
            .I(N__32030));
    LocalMux I__5924 (
            .O(N__32030),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__5923 (
            .O(N__32027),
            .I(N__32024));
    InMux I__5922 (
            .O(N__32024),
            .I(N__32021));
    LocalMux I__5921 (
            .O(N__32021),
            .I(N__32018));
    Span4Mux_h I__5920 (
            .O(N__32018),
            .I(N__32015));
    Odrv4 I__5919 (
            .O(N__32015),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ1Z_6 ));
    InMux I__5918 (
            .O(N__32012),
            .I(N__32008));
    InMux I__5917 (
            .O(N__32011),
            .I(N__32005));
    LocalMux I__5916 (
            .O(N__32008),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__5915 (
            .O(N__32005),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__5914 (
            .O(N__32000),
            .I(N__31997));
    LocalMux I__5913 (
            .O(N__31997),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__5912 (
            .O(N__31994),
            .I(N__31990));
    InMux I__5911 (
            .O(N__31993),
            .I(N__31987));
    LocalMux I__5910 (
            .O(N__31990),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__5909 (
            .O(N__31987),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__5908 (
            .O(N__31982),
            .I(N__31979));
    LocalMux I__5907 (
            .O(N__31979),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__5906 (
            .O(N__31976),
            .I(N__31973));
    LocalMux I__5905 (
            .O(N__31973),
            .I(N__31969));
    InMux I__5904 (
            .O(N__31972),
            .I(N__31966));
    Odrv4 I__5903 (
            .O(N__31969),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__5902 (
            .O(N__31966),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__5901 (
            .O(N__31961),
            .I(N__31958));
    LocalMux I__5900 (
            .O(N__31958),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__5899 (
            .O(N__31955),
            .I(N__31952));
    InMux I__5898 (
            .O(N__31952),
            .I(N__31949));
    LocalMux I__5897 (
            .O(N__31949),
            .I(N__31946));
    Span4Mux_h I__5896 (
            .O(N__31946),
            .I(N__31943));
    Odrv4 I__5895 (
            .O(N__31943),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__5894 (
            .O(N__31940),
            .I(N__31937));
    LocalMux I__5893 (
            .O(N__31937),
            .I(N__31933));
    InMux I__5892 (
            .O(N__31936),
            .I(N__31930));
    Odrv4 I__5891 (
            .O(N__31933),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__5890 (
            .O(N__31930),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__5889 (
            .O(N__31925),
            .I(N__31922));
    LocalMux I__5888 (
            .O(N__31922),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__5887 (
            .O(N__31919),
            .I(N__31913));
    InMux I__5886 (
            .O(N__31918),
            .I(N__31909));
    InMux I__5885 (
            .O(N__31917),
            .I(N__31906));
    CascadeMux I__5884 (
            .O(N__31916),
            .I(N__31903));
    LocalMux I__5883 (
            .O(N__31913),
            .I(N__31900));
    InMux I__5882 (
            .O(N__31912),
            .I(N__31897));
    LocalMux I__5881 (
            .O(N__31909),
            .I(N__31894));
    LocalMux I__5880 (
            .O(N__31906),
            .I(N__31891));
    InMux I__5879 (
            .O(N__31903),
            .I(N__31888));
    Span4Mux_v I__5878 (
            .O(N__31900),
            .I(N__31885));
    LocalMux I__5877 (
            .O(N__31897),
            .I(N__31882));
    Span4Mux_v I__5876 (
            .O(N__31894),
            .I(N__31877));
    Span4Mux_v I__5875 (
            .O(N__31891),
            .I(N__31877));
    LocalMux I__5874 (
            .O(N__31888),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__5873 (
            .O(N__31885),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__5872 (
            .O(N__31882),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__5871 (
            .O(N__31877),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__5870 (
            .O(N__31868),
            .I(N__31865));
    InMux I__5869 (
            .O(N__31865),
            .I(N__31862));
    LocalMux I__5868 (
            .O(N__31862),
            .I(N__31859));
    Odrv4 I__5867 (
            .O(N__31859),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    CascadeMux I__5866 (
            .O(N__31856),
            .I(N__31851));
    CascadeMux I__5865 (
            .O(N__31855),
            .I(N__31848));
    InMux I__5864 (
            .O(N__31854),
            .I(N__31843));
    InMux I__5863 (
            .O(N__31851),
            .I(N__31840));
    InMux I__5862 (
            .O(N__31848),
            .I(N__31837));
    InMux I__5861 (
            .O(N__31847),
            .I(N__31834));
    InMux I__5860 (
            .O(N__31846),
            .I(N__31831));
    LocalMux I__5859 (
            .O(N__31843),
            .I(N__31828));
    LocalMux I__5858 (
            .O(N__31840),
            .I(N__31825));
    LocalMux I__5857 (
            .O(N__31837),
            .I(N__31822));
    LocalMux I__5856 (
            .O(N__31834),
            .I(N__31819));
    LocalMux I__5855 (
            .O(N__31831),
            .I(N__31814));
    Span4Mux_h I__5854 (
            .O(N__31828),
            .I(N__31814));
    Span4Mux_h I__5853 (
            .O(N__31825),
            .I(N__31809));
    Span4Mux_v I__5852 (
            .O(N__31822),
            .I(N__31809));
    Span4Mux_h I__5851 (
            .O(N__31819),
            .I(N__31806));
    Span4Mux_v I__5850 (
            .O(N__31814),
            .I(N__31803));
    Odrv4 I__5849 (
            .O(N__31809),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__5848 (
            .O(N__31806),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__5847 (
            .O(N__31803),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    CascadeMux I__5846 (
            .O(N__31796),
            .I(N__31792));
    InMux I__5845 (
            .O(N__31795),
            .I(N__31789));
    InMux I__5844 (
            .O(N__31792),
            .I(N__31786));
    LocalMux I__5843 (
            .O(N__31789),
            .I(N__31781));
    LocalMux I__5842 (
            .O(N__31786),
            .I(N__31778));
    CascadeMux I__5841 (
            .O(N__31785),
            .I(N__31775));
    InMux I__5840 (
            .O(N__31784),
            .I(N__31771));
    Span4Mux_v I__5839 (
            .O(N__31781),
            .I(N__31768));
    Span4Mux_v I__5838 (
            .O(N__31778),
            .I(N__31765));
    InMux I__5837 (
            .O(N__31775),
            .I(N__31762));
    InMux I__5836 (
            .O(N__31774),
            .I(N__31759));
    LocalMux I__5835 (
            .O(N__31771),
            .I(N__31756));
    Odrv4 I__5834 (
            .O(N__31768),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__5833 (
            .O(N__31765),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__5832 (
            .O(N__31762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__5831 (
            .O(N__31759),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__5830 (
            .O(N__31756),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__5829 (
            .O(N__31745),
            .I(N__31741));
    CascadeMux I__5828 (
            .O(N__31744),
            .I(N__31736));
    InMux I__5827 (
            .O(N__31741),
            .I(N__31732));
    InMux I__5826 (
            .O(N__31740),
            .I(N__31729));
    InMux I__5825 (
            .O(N__31739),
            .I(N__31726));
    InMux I__5824 (
            .O(N__31736),
            .I(N__31723));
    InMux I__5823 (
            .O(N__31735),
            .I(N__31720));
    LocalMux I__5822 (
            .O(N__31732),
            .I(N__31717));
    LocalMux I__5821 (
            .O(N__31729),
            .I(N__31714));
    LocalMux I__5820 (
            .O(N__31726),
            .I(N__31711));
    LocalMux I__5819 (
            .O(N__31723),
            .I(N__31708));
    LocalMux I__5818 (
            .O(N__31720),
            .I(N__31705));
    Span4Mux_v I__5817 (
            .O(N__31717),
            .I(N__31702));
    Span4Mux_h I__5816 (
            .O(N__31714),
            .I(N__31697));
    Span4Mux_h I__5815 (
            .O(N__31711),
            .I(N__31697));
    Span4Mux_h I__5814 (
            .O(N__31708),
            .I(N__31692));
    Span4Mux_v I__5813 (
            .O(N__31705),
            .I(N__31692));
    Odrv4 I__5812 (
            .O(N__31702),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__5811 (
            .O(N__31697),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__5810 (
            .O(N__31692),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__5809 (
            .O(N__31685),
            .I(N__31679));
    CascadeMux I__5808 (
            .O(N__31684),
            .I(N__31675));
    InMux I__5807 (
            .O(N__31683),
            .I(N__31670));
    InMux I__5806 (
            .O(N__31682),
            .I(N__31670));
    LocalMux I__5805 (
            .O(N__31679),
            .I(N__31667));
    InMux I__5804 (
            .O(N__31678),
            .I(N__31664));
    InMux I__5803 (
            .O(N__31675),
            .I(N__31661));
    LocalMux I__5802 (
            .O(N__31670),
            .I(N__31658));
    Span4Mux_v I__5801 (
            .O(N__31667),
            .I(N__31655));
    LocalMux I__5800 (
            .O(N__31664),
            .I(N__31652));
    LocalMux I__5799 (
            .O(N__31661),
            .I(N__31647));
    Span4Mux_v I__5798 (
            .O(N__31658),
            .I(N__31647));
    Odrv4 I__5797 (
            .O(N__31655),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5796 (
            .O(N__31652),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5795 (
            .O(N__31647),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__5794 (
            .O(N__31640),
            .I(N__31637));
    LocalMux I__5793 (
            .O(N__31637),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    InMux I__5792 (
            .O(N__31634),
            .I(N__31631));
    LocalMux I__5791 (
            .O(N__31631),
            .I(N__31627));
    InMux I__5790 (
            .O(N__31630),
            .I(N__31624));
    Span4Mux_h I__5789 (
            .O(N__31627),
            .I(N__31621));
    LocalMux I__5788 (
            .O(N__31624),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__5787 (
            .O(N__31621),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    CascadeMux I__5786 (
            .O(N__31616),
            .I(N__31612));
    InMux I__5785 (
            .O(N__31615),
            .I(N__31608));
    InMux I__5784 (
            .O(N__31612),
            .I(N__31605));
    InMux I__5783 (
            .O(N__31611),
            .I(N__31602));
    LocalMux I__5782 (
            .O(N__31608),
            .I(N__31597));
    LocalMux I__5781 (
            .O(N__31605),
            .I(N__31592));
    LocalMux I__5780 (
            .O(N__31602),
            .I(N__31592));
    InMux I__5779 (
            .O(N__31601),
            .I(N__31587));
    InMux I__5778 (
            .O(N__31600),
            .I(N__31587));
    Span12Mux_v I__5777 (
            .O(N__31597),
            .I(N__31584));
    Span4Mux_h I__5776 (
            .O(N__31592),
            .I(N__31581));
    LocalMux I__5775 (
            .O(N__31587),
            .I(N__31578));
    Odrv12 I__5774 (
            .O(N__31584),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5773 (
            .O(N__31581),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5772 (
            .O(N__31578),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__5771 (
            .O(N__31571),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16_cascade_ ));
    InMux I__5770 (
            .O(N__31568),
            .I(N__31565));
    LocalMux I__5769 (
            .O(N__31565),
            .I(N__31562));
    Span4Mux_h I__5768 (
            .O(N__31562),
            .I(N__31559));
    Odrv4 I__5767 (
            .O(N__31559),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__5766 (
            .O(N__31556),
            .I(N__31553));
    LocalMux I__5765 (
            .O(N__31553),
            .I(N__31550));
    Odrv4 I__5764 (
            .O(N__31550),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ));
    InMux I__5763 (
            .O(N__31547),
            .I(N__31543));
    InMux I__5762 (
            .O(N__31546),
            .I(N__31540));
    LocalMux I__5761 (
            .O(N__31543),
            .I(N__31534));
    LocalMux I__5760 (
            .O(N__31540),
            .I(N__31534));
    InMux I__5759 (
            .O(N__31539),
            .I(N__31531));
    Span4Mux_h I__5758 (
            .O(N__31534),
            .I(N__31528));
    LocalMux I__5757 (
            .O(N__31531),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv4 I__5756 (
            .O(N__31528),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    InMux I__5755 (
            .O(N__31523),
            .I(N__31494));
    InMux I__5754 (
            .O(N__31522),
            .I(N__31489));
    InMux I__5753 (
            .O(N__31521),
            .I(N__31489));
    InMux I__5752 (
            .O(N__31520),
            .I(N__31482));
    InMux I__5751 (
            .O(N__31519),
            .I(N__31482));
    InMux I__5750 (
            .O(N__31518),
            .I(N__31482));
    InMux I__5749 (
            .O(N__31517),
            .I(N__31479));
    InMux I__5748 (
            .O(N__31516),
            .I(N__31470));
    InMux I__5747 (
            .O(N__31515),
            .I(N__31470));
    InMux I__5746 (
            .O(N__31514),
            .I(N__31470));
    InMux I__5745 (
            .O(N__31513),
            .I(N__31470));
    InMux I__5744 (
            .O(N__31512),
            .I(N__31466));
    InMux I__5743 (
            .O(N__31511),
            .I(N__31463));
    InMux I__5742 (
            .O(N__31510),
            .I(N__31448));
    InMux I__5741 (
            .O(N__31509),
            .I(N__31448));
    InMux I__5740 (
            .O(N__31508),
            .I(N__31448));
    InMux I__5739 (
            .O(N__31507),
            .I(N__31448));
    InMux I__5738 (
            .O(N__31506),
            .I(N__31448));
    InMux I__5737 (
            .O(N__31505),
            .I(N__31448));
    InMux I__5736 (
            .O(N__31504),
            .I(N__31448));
    InMux I__5735 (
            .O(N__31503),
            .I(N__31433));
    InMux I__5734 (
            .O(N__31502),
            .I(N__31433));
    InMux I__5733 (
            .O(N__31501),
            .I(N__31433));
    InMux I__5732 (
            .O(N__31500),
            .I(N__31433));
    InMux I__5731 (
            .O(N__31499),
            .I(N__31433));
    InMux I__5730 (
            .O(N__31498),
            .I(N__31433));
    InMux I__5729 (
            .O(N__31497),
            .I(N__31433));
    LocalMux I__5728 (
            .O(N__31494),
            .I(N__31418));
    LocalMux I__5727 (
            .O(N__31489),
            .I(N__31415));
    LocalMux I__5726 (
            .O(N__31482),
            .I(N__31408));
    LocalMux I__5725 (
            .O(N__31479),
            .I(N__31408));
    LocalMux I__5724 (
            .O(N__31470),
            .I(N__31408));
    InMux I__5723 (
            .O(N__31469),
            .I(N__31405));
    LocalMux I__5722 (
            .O(N__31466),
            .I(N__31402));
    LocalMux I__5721 (
            .O(N__31463),
            .I(N__31384));
    LocalMux I__5720 (
            .O(N__31448),
            .I(N__31384));
    LocalMux I__5719 (
            .O(N__31433),
            .I(N__31384));
    InMux I__5718 (
            .O(N__31432),
            .I(N__31375));
    InMux I__5717 (
            .O(N__31431),
            .I(N__31375));
    InMux I__5716 (
            .O(N__31430),
            .I(N__31375));
    InMux I__5715 (
            .O(N__31429),
            .I(N__31375));
    InMux I__5714 (
            .O(N__31428),
            .I(N__31372));
    InMux I__5713 (
            .O(N__31427),
            .I(N__31357));
    InMux I__5712 (
            .O(N__31426),
            .I(N__31357));
    InMux I__5711 (
            .O(N__31425),
            .I(N__31357));
    InMux I__5710 (
            .O(N__31424),
            .I(N__31357));
    InMux I__5709 (
            .O(N__31423),
            .I(N__31357));
    InMux I__5708 (
            .O(N__31422),
            .I(N__31357));
    InMux I__5707 (
            .O(N__31421),
            .I(N__31357));
    Span4Mux_v I__5706 (
            .O(N__31418),
            .I(N__31352));
    Span4Mux_v I__5705 (
            .O(N__31415),
            .I(N__31352));
    Span4Mux_h I__5704 (
            .O(N__31408),
            .I(N__31349));
    LocalMux I__5703 (
            .O(N__31405),
            .I(N__31344));
    Span4Mux_v I__5702 (
            .O(N__31402),
            .I(N__31344));
    InMux I__5701 (
            .O(N__31401),
            .I(N__31329));
    InMux I__5700 (
            .O(N__31400),
            .I(N__31329));
    InMux I__5699 (
            .O(N__31399),
            .I(N__31329));
    InMux I__5698 (
            .O(N__31398),
            .I(N__31329));
    InMux I__5697 (
            .O(N__31397),
            .I(N__31329));
    InMux I__5696 (
            .O(N__31396),
            .I(N__31329));
    InMux I__5695 (
            .O(N__31395),
            .I(N__31329));
    InMux I__5694 (
            .O(N__31394),
            .I(N__31320));
    InMux I__5693 (
            .O(N__31393),
            .I(N__31320));
    InMux I__5692 (
            .O(N__31392),
            .I(N__31320));
    InMux I__5691 (
            .O(N__31391),
            .I(N__31320));
    Span4Mux_v I__5690 (
            .O(N__31384),
            .I(N__31315));
    LocalMux I__5689 (
            .O(N__31375),
            .I(N__31315));
    LocalMux I__5688 (
            .O(N__31372),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    LocalMux I__5687 (
            .O(N__31357),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__5686 (
            .O(N__31352),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__5685 (
            .O(N__31349),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__5684 (
            .O(N__31344),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    LocalMux I__5683 (
            .O(N__31329),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    LocalMux I__5682 (
            .O(N__31320),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__5681 (
            .O(N__31315),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__5680 (
            .O(N__31298),
            .I(N__31295));
    LocalMux I__5679 (
            .O(N__31295),
            .I(N__31290));
    InMux I__5678 (
            .O(N__31294),
            .I(N__31287));
    InMux I__5677 (
            .O(N__31293),
            .I(N__31284));
    Span4Mux_h I__5676 (
            .O(N__31290),
            .I(N__31281));
    LocalMux I__5675 (
            .O(N__31287),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    LocalMux I__5674 (
            .O(N__31284),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv4 I__5673 (
            .O(N__31281),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    InMux I__5672 (
            .O(N__31274),
            .I(N__31271));
    LocalMux I__5671 (
            .O(N__31271),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__5670 (
            .O(N__31268),
            .I(N__31264));
    InMux I__5669 (
            .O(N__31267),
            .I(N__31261));
    InMux I__5668 (
            .O(N__31264),
            .I(N__31257));
    LocalMux I__5667 (
            .O(N__31261),
            .I(N__31254));
    InMux I__5666 (
            .O(N__31260),
            .I(N__31251));
    LocalMux I__5665 (
            .O(N__31257),
            .I(N__31246));
    Span4Mux_h I__5664 (
            .O(N__31254),
            .I(N__31243));
    LocalMux I__5663 (
            .O(N__31251),
            .I(N__31240));
    InMux I__5662 (
            .O(N__31250),
            .I(N__31235));
    InMux I__5661 (
            .O(N__31249),
            .I(N__31235));
    Odrv12 I__5660 (
            .O(N__31246),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__5659 (
            .O(N__31243),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__5658 (
            .O(N__31240),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__5657 (
            .O(N__31235),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__5656 (
            .O(N__31226),
            .I(N__31223));
    LocalMux I__5655 (
            .O(N__31223),
            .I(N__31220));
    Odrv4 I__5654 (
            .O(N__31220),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    InMux I__5653 (
            .O(N__31217),
            .I(N__31214));
    LocalMux I__5652 (
            .O(N__31214),
            .I(N__31211));
    Span4Mux_h I__5651 (
            .O(N__31211),
            .I(N__31208));
    Odrv4 I__5650 (
            .O(N__31208),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ));
    InMux I__5649 (
            .O(N__31205),
            .I(N__31201));
    InMux I__5648 (
            .O(N__31204),
            .I(N__31198));
    LocalMux I__5647 (
            .O(N__31201),
            .I(N__31195));
    LocalMux I__5646 (
            .O(N__31198),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    Odrv4 I__5645 (
            .O(N__31195),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    InMux I__5644 (
            .O(N__31190),
            .I(N__31186));
    InMux I__5643 (
            .O(N__31189),
            .I(N__31182));
    LocalMux I__5642 (
            .O(N__31186),
            .I(N__31178));
    InMux I__5641 (
            .O(N__31185),
            .I(N__31174));
    LocalMux I__5640 (
            .O(N__31182),
            .I(N__31171));
    InMux I__5639 (
            .O(N__31181),
            .I(N__31168));
    Span4Mux_h I__5638 (
            .O(N__31178),
            .I(N__31165));
    InMux I__5637 (
            .O(N__31177),
            .I(N__31162));
    LocalMux I__5636 (
            .O(N__31174),
            .I(N__31159));
    Span12Mux_v I__5635 (
            .O(N__31171),
            .I(N__31154));
    LocalMux I__5634 (
            .O(N__31168),
            .I(N__31154));
    Odrv4 I__5633 (
            .O(N__31165),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__5632 (
            .O(N__31162),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__5631 (
            .O(N__31159),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv12 I__5630 (
            .O(N__31154),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__5629 (
            .O(N__31145),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18_cascade_ ));
    InMux I__5628 (
            .O(N__31142),
            .I(N__31139));
    LocalMux I__5627 (
            .O(N__31139),
            .I(N__31136));
    Odrv4 I__5626 (
            .O(N__31136),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__5625 (
            .O(N__31133),
            .I(N__31130));
    LocalMux I__5624 (
            .O(N__31130),
            .I(N__31127));
    Span4Mux_h I__5623 (
            .O(N__31127),
            .I(N__31124));
    Odrv4 I__5622 (
            .O(N__31124),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ));
    InMux I__5621 (
            .O(N__31121),
            .I(N__31118));
    LocalMux I__5620 (
            .O(N__31118),
            .I(N__31113));
    InMux I__5619 (
            .O(N__31117),
            .I(N__31110));
    InMux I__5618 (
            .O(N__31116),
            .I(N__31107));
    Span4Mux_v I__5617 (
            .O(N__31113),
            .I(N__31104));
    LocalMux I__5616 (
            .O(N__31110),
            .I(N__31101));
    LocalMux I__5615 (
            .O(N__31107),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__5614 (
            .O(N__31104),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__5613 (
            .O(N__31101),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    InMux I__5612 (
            .O(N__31094),
            .I(N__31090));
    InMux I__5611 (
            .O(N__31093),
            .I(N__31087));
    LocalMux I__5610 (
            .O(N__31090),
            .I(N__31081));
    LocalMux I__5609 (
            .O(N__31087),
            .I(N__31081));
    InMux I__5608 (
            .O(N__31086),
            .I(N__31078));
    Span4Mux_v I__5607 (
            .O(N__31081),
            .I(N__31075));
    LocalMux I__5606 (
            .O(N__31078),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    Odrv4 I__5605 (
            .O(N__31075),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    InMux I__5604 (
            .O(N__31070),
            .I(N__31067));
    LocalMux I__5603 (
            .O(N__31067),
            .I(N__31064));
    Span4Mux_v I__5602 (
            .O(N__31064),
            .I(N__31059));
    InMux I__5601 (
            .O(N__31063),
            .I(N__31056));
    InMux I__5600 (
            .O(N__31062),
            .I(N__31053));
    Span4Mux_v I__5599 (
            .O(N__31059),
            .I(N__31048));
    LocalMux I__5598 (
            .O(N__31056),
            .I(N__31048));
    LocalMux I__5597 (
            .O(N__31053),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv4 I__5596 (
            .O(N__31048),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    InMux I__5595 (
            .O(N__31043),
            .I(N__31039));
    InMux I__5594 (
            .O(N__31042),
            .I(N__31036));
    LocalMux I__5593 (
            .O(N__31039),
            .I(N__31032));
    LocalMux I__5592 (
            .O(N__31036),
            .I(N__31029));
    InMux I__5591 (
            .O(N__31035),
            .I(N__31026));
    Span4Mux_h I__5590 (
            .O(N__31032),
            .I(N__31023));
    Span4Mux_h I__5589 (
            .O(N__31029),
            .I(N__31020));
    LocalMux I__5588 (
            .O(N__31026),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__5587 (
            .O(N__31023),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__5586 (
            .O(N__31020),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__5585 (
            .O(N__31013),
            .I(N__31010));
    LocalMux I__5584 (
            .O(N__31010),
            .I(N__31007));
    Span4Mux_v I__5583 (
            .O(N__31007),
            .I(N__31004));
    Odrv4 I__5582 (
            .O(N__31004),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    CascadeMux I__5581 (
            .O(N__31001),
            .I(N__30998));
    InMux I__5580 (
            .O(N__30998),
            .I(N__30995));
    LocalMux I__5579 (
            .O(N__30995),
            .I(N__30992));
    Span4Mux_v I__5578 (
            .O(N__30992),
            .I(N__30989));
    Odrv4 I__5577 (
            .O(N__30989),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__5576 (
            .O(N__30986),
            .I(N__30983));
    LocalMux I__5575 (
            .O(N__30983),
            .I(N__30980));
    Span4Mux_h I__5574 (
            .O(N__30980),
            .I(N__30977));
    Span4Mux_h I__5573 (
            .O(N__30977),
            .I(N__30974));
    Odrv4 I__5572 (
            .O(N__30974),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ));
    CascadeMux I__5571 (
            .O(N__30971),
            .I(N__30968));
    InMux I__5570 (
            .O(N__30968),
            .I(N__30965));
    LocalMux I__5569 (
            .O(N__30965),
            .I(N__30962));
    Span4Mux_h I__5568 (
            .O(N__30962),
            .I(N__30959));
    Span4Mux_h I__5567 (
            .O(N__30959),
            .I(N__30956));
    Odrv4 I__5566 (
            .O(N__30956),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__5565 (
            .O(N__30953),
            .I(N__30950));
    InMux I__5564 (
            .O(N__30950),
            .I(N__30947));
    LocalMux I__5563 (
            .O(N__30947),
            .I(N__30944));
    Span4Mux_h I__5562 (
            .O(N__30944),
            .I(N__30941));
    Odrv4 I__5561 (
            .O(N__30941),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    InMux I__5560 (
            .O(N__30938),
            .I(N__30928));
    InMux I__5559 (
            .O(N__30937),
            .I(N__30928));
    InMux I__5558 (
            .O(N__30936),
            .I(N__30924));
    InMux I__5557 (
            .O(N__30935),
            .I(N__30917));
    InMux I__5556 (
            .O(N__30934),
            .I(N__30917));
    InMux I__5555 (
            .O(N__30933),
            .I(N__30917));
    LocalMux I__5554 (
            .O(N__30928),
            .I(N__30914));
    InMux I__5553 (
            .O(N__30927),
            .I(N__30911));
    LocalMux I__5552 (
            .O(N__30924),
            .I(\delay_measurement_inst.N_299 ));
    LocalMux I__5551 (
            .O(N__30917),
            .I(\delay_measurement_inst.N_299 ));
    Odrv4 I__5550 (
            .O(N__30914),
            .I(\delay_measurement_inst.N_299 ));
    LocalMux I__5549 (
            .O(N__30911),
            .I(\delay_measurement_inst.N_299 ));
    CascadeMux I__5548 (
            .O(N__30902),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_ ));
    InMux I__5547 (
            .O(N__30899),
            .I(N__30896));
    LocalMux I__5546 (
            .O(N__30896),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ));
    CascadeMux I__5545 (
            .O(N__30893),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9_cascade_ ));
    CascadeMux I__5544 (
            .O(N__30890),
            .I(N__30886));
    CascadeMux I__5543 (
            .O(N__30889),
            .I(N__30883));
    InMux I__5542 (
            .O(N__30886),
            .I(N__30880));
    InMux I__5541 (
            .O(N__30883),
            .I(N__30877));
    LocalMux I__5540 (
            .O(N__30880),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ));
    LocalMux I__5539 (
            .O(N__30877),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ));
    CEMux I__5538 (
            .O(N__30872),
            .I(N__30865));
    CEMux I__5537 (
            .O(N__30871),
            .I(N__30862));
    CEMux I__5536 (
            .O(N__30870),
            .I(N__30859));
    CEMux I__5535 (
            .O(N__30869),
            .I(N__30856));
    CEMux I__5534 (
            .O(N__30868),
            .I(N__30853));
    LocalMux I__5533 (
            .O(N__30865),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__5532 (
            .O(N__30862),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__5531 (
            .O(N__30859),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__5530 (
            .O(N__30856),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__5529 (
            .O(N__30853),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    CascadeMux I__5528 (
            .O(N__30842),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_ ));
    InMux I__5527 (
            .O(N__30839),
            .I(N__30836));
    LocalMux I__5526 (
            .O(N__30836),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ));
    InMux I__5525 (
            .O(N__30833),
            .I(N__30830));
    LocalMux I__5524 (
            .O(N__30830),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ));
    InMux I__5523 (
            .O(N__30827),
            .I(N__30824));
    LocalMux I__5522 (
            .O(N__30824),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7 ));
    InMux I__5521 (
            .O(N__30821),
            .I(N__30818));
    LocalMux I__5520 (
            .O(N__30818),
            .I(N__30815));
    Span4Mux_h I__5519 (
            .O(N__30815),
            .I(N__30812));
    Odrv4 I__5518 (
            .O(N__30812),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ));
    CascadeMux I__5517 (
            .O(N__30809),
            .I(N__30806));
    InMux I__5516 (
            .O(N__30806),
            .I(N__30803));
    LocalMux I__5515 (
            .O(N__30803),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ));
    InMux I__5514 (
            .O(N__30800),
            .I(N__30797));
    LocalMux I__5513 (
            .O(N__30797),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    CascadeMux I__5512 (
            .O(N__30794),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ));
    InMux I__5511 (
            .O(N__30791),
            .I(N__30788));
    LocalMux I__5510 (
            .O(N__30788),
            .I(N__30785));
    Odrv4 I__5509 (
            .O(N__30785),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ));
    CascadeMux I__5508 (
            .O(N__30782),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ));
    CascadeMux I__5507 (
            .O(N__30779),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6_cascade_ ));
    InMux I__5506 (
            .O(N__30776),
            .I(N__30773));
    LocalMux I__5505 (
            .O(N__30773),
            .I(\delay_measurement_inst.N_42 ));
    InMux I__5504 (
            .O(N__30770),
            .I(N__30767));
    LocalMux I__5503 (
            .O(N__30767),
            .I(N__30761));
    InMux I__5502 (
            .O(N__30766),
            .I(N__30758));
    InMux I__5501 (
            .O(N__30765),
            .I(N__30755));
    CascadeMux I__5500 (
            .O(N__30764),
            .I(N__30752));
    Span4Mux_h I__5499 (
            .O(N__30761),
            .I(N__30749));
    LocalMux I__5498 (
            .O(N__30758),
            .I(N__30743));
    LocalMux I__5497 (
            .O(N__30755),
            .I(N__30743));
    InMux I__5496 (
            .O(N__30752),
            .I(N__30740));
    Span4Mux_h I__5495 (
            .O(N__30749),
            .I(N__30737));
    InMux I__5494 (
            .O(N__30748),
            .I(N__30734));
    Span4Mux_h I__5493 (
            .O(N__30743),
            .I(N__30731));
    LocalMux I__5492 (
            .O(N__30740),
            .I(N__30728));
    Odrv4 I__5491 (
            .O(N__30737),
            .I(measured_delay_hc_18));
    LocalMux I__5490 (
            .O(N__30734),
            .I(measured_delay_hc_18));
    Odrv4 I__5489 (
            .O(N__30731),
            .I(measured_delay_hc_18));
    Odrv4 I__5488 (
            .O(N__30728),
            .I(measured_delay_hc_18));
    InMux I__5487 (
            .O(N__30719),
            .I(N__30716));
    LocalMux I__5486 (
            .O(N__30716),
            .I(\delay_measurement_inst.N_26 ));
    InMux I__5485 (
            .O(N__30713),
            .I(N__30710));
    LocalMux I__5484 (
            .O(N__30710),
            .I(N__30707));
    Span4Mux_h I__5483 (
            .O(N__30707),
            .I(N__30704));
    Span4Mux_v I__5482 (
            .O(N__30704),
            .I(N__30699));
    InMux I__5481 (
            .O(N__30703),
            .I(N__30696));
    InMux I__5480 (
            .O(N__30702),
            .I(N__30693));
    Odrv4 I__5479 (
            .O(N__30699),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__5478 (
            .O(N__30696),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__5477 (
            .O(N__30693),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__5476 (
            .O(N__30686),
            .I(N__30683));
    LocalMux I__5475 (
            .O(N__30683),
            .I(N__30680));
    Span4Mux_v I__5474 (
            .O(N__30680),
            .I(N__30674));
    InMux I__5473 (
            .O(N__30679),
            .I(N__30669));
    InMux I__5472 (
            .O(N__30678),
            .I(N__30669));
    InMux I__5471 (
            .O(N__30677),
            .I(N__30666));
    Odrv4 I__5470 (
            .O(N__30674),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5469 (
            .O(N__30669),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5468 (
            .O(N__30666),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__5467 (
            .O(N__30659),
            .I(N__30656));
    LocalMux I__5466 (
            .O(N__30656),
            .I(N__30653));
    Span4Mux_h I__5465 (
            .O(N__30653),
            .I(N__30650));
    Odrv4 I__5464 (
            .O(N__30650),
            .I(\delay_measurement_inst.N_27 ));
    InMux I__5463 (
            .O(N__30647),
            .I(N__30644));
    LocalMux I__5462 (
            .O(N__30644),
            .I(N__30641));
    Span4Mux_h I__5461 (
            .O(N__30641),
            .I(N__30637));
    InMux I__5460 (
            .O(N__30640),
            .I(N__30634));
    Odrv4 I__5459 (
            .O(N__30637),
            .I(\delay_measurement_inst.elapsed_time_hc_29 ));
    LocalMux I__5458 (
            .O(N__30634),
            .I(\delay_measurement_inst.elapsed_time_hc_29 ));
    InMux I__5457 (
            .O(N__30629),
            .I(N__30626));
    LocalMux I__5456 (
            .O(N__30626),
            .I(\delay_measurement_inst.N_53 ));
    InMux I__5455 (
            .O(N__30623),
            .I(N__30619));
    InMux I__5454 (
            .O(N__30622),
            .I(N__30616));
    LocalMux I__5453 (
            .O(N__30619),
            .I(measured_delay_hc_29));
    LocalMux I__5452 (
            .O(N__30616),
            .I(measured_delay_hc_29));
    InMux I__5451 (
            .O(N__30611),
            .I(N__30608));
    LocalMux I__5450 (
            .O(N__30608),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3 ));
    InMux I__5449 (
            .O(N__30605),
            .I(N__30602));
    LocalMux I__5448 (
            .O(N__30602),
            .I(\delay_measurement_inst.N_54 ));
    InMux I__5447 (
            .O(N__30599),
            .I(N__30595));
    InMux I__5446 (
            .O(N__30598),
            .I(N__30592));
    LocalMux I__5445 (
            .O(N__30595),
            .I(measured_delay_hc_30));
    LocalMux I__5444 (
            .O(N__30592),
            .I(measured_delay_hc_30));
    InMux I__5443 (
            .O(N__30587),
            .I(N__30584));
    LocalMux I__5442 (
            .O(N__30584),
            .I(N__30581));
    Span4Mux_h I__5441 (
            .O(N__30581),
            .I(N__30578));
    Odrv4 I__5440 (
            .O(N__30578),
            .I(delay_hc_input_c));
    InMux I__5439 (
            .O(N__30575),
            .I(N__30572));
    LocalMux I__5438 (
            .O(N__30572),
            .I(delay_hc_d1));
    InMux I__5437 (
            .O(N__30569),
            .I(N__30566));
    LocalMux I__5436 (
            .O(N__30566),
            .I(N__30560));
    InMux I__5435 (
            .O(N__30565),
            .I(N__30555));
    InMux I__5434 (
            .O(N__30564),
            .I(N__30555));
    InMux I__5433 (
            .O(N__30563),
            .I(N__30552));
    Span4Mux_h I__5432 (
            .O(N__30560),
            .I(N__30547));
    LocalMux I__5431 (
            .O(N__30555),
            .I(N__30547));
    LocalMux I__5430 (
            .O(N__30552),
            .I(N__30544));
    Span4Mux_v I__5429 (
            .O(N__30547),
            .I(N__30541));
    Span4Mux_h I__5428 (
            .O(N__30544),
            .I(N__30538));
    Odrv4 I__5427 (
            .O(N__30541),
            .I(delay_hc_d2));
    Odrv4 I__5426 (
            .O(N__30538),
            .I(delay_hc_d2));
    InMux I__5425 (
            .O(N__30533),
            .I(N__30530));
    LocalMux I__5424 (
            .O(N__30530),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ));
    CascadeMux I__5423 (
            .O(N__30527),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_ ));
    InMux I__5422 (
            .O(N__30524),
            .I(N__30521));
    LocalMux I__5421 (
            .O(N__30521),
            .I(N__30518));
    Odrv4 I__5420 (
            .O(N__30518),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ));
    InMux I__5419 (
            .O(N__30515),
            .I(N__30512));
    LocalMux I__5418 (
            .O(N__30512),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3 ));
    CascadeMux I__5417 (
            .O(N__30509),
            .I(N__30506));
    InMux I__5416 (
            .O(N__30506),
            .I(N__30501));
    InMux I__5415 (
            .O(N__30505),
            .I(N__30498));
    InMux I__5414 (
            .O(N__30504),
            .I(N__30495));
    LocalMux I__5413 (
            .O(N__30501),
            .I(measured_delay_hc_20));
    LocalMux I__5412 (
            .O(N__30498),
            .I(measured_delay_hc_20));
    LocalMux I__5411 (
            .O(N__30495),
            .I(measured_delay_hc_20));
    InMux I__5410 (
            .O(N__30488),
            .I(N__30483));
    InMux I__5409 (
            .O(N__30487),
            .I(N__30480));
    CascadeMux I__5408 (
            .O(N__30486),
            .I(N__30477));
    LocalMux I__5407 (
            .O(N__30483),
            .I(N__30474));
    LocalMux I__5406 (
            .O(N__30480),
            .I(N__30471));
    InMux I__5405 (
            .O(N__30477),
            .I(N__30468));
    Span4Mux_h I__5404 (
            .O(N__30474),
            .I(N__30463));
    Span4Mux_v I__5403 (
            .O(N__30471),
            .I(N__30463));
    LocalMux I__5402 (
            .O(N__30468),
            .I(N__30460));
    Odrv4 I__5401 (
            .O(N__30463),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    Odrv4 I__5400 (
            .O(N__30460),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    CascadeMux I__5399 (
            .O(N__30455),
            .I(\delay_measurement_inst.N_29_cascade_ ));
    CascadeMux I__5398 (
            .O(N__30452),
            .I(N__30448));
    CascadeMux I__5397 (
            .O(N__30451),
            .I(N__30444));
    InMux I__5396 (
            .O(N__30448),
            .I(N__30441));
    InMux I__5395 (
            .O(N__30447),
            .I(N__30438));
    InMux I__5394 (
            .O(N__30444),
            .I(N__30435));
    LocalMux I__5393 (
            .O(N__30441),
            .I(N__30431));
    LocalMux I__5392 (
            .O(N__30438),
            .I(N__30426));
    LocalMux I__5391 (
            .O(N__30435),
            .I(N__30426));
    InMux I__5390 (
            .O(N__30434),
            .I(N__30423));
    Span4Mux_v I__5389 (
            .O(N__30431),
            .I(N__30419));
    Span4Mux_v I__5388 (
            .O(N__30426),
            .I(N__30414));
    LocalMux I__5387 (
            .O(N__30423),
            .I(N__30414));
    InMux I__5386 (
            .O(N__30422),
            .I(N__30411));
    Span4Mux_v I__5385 (
            .O(N__30419),
            .I(N__30408));
    Span4Mux_v I__5384 (
            .O(N__30414),
            .I(N__30405));
    LocalMux I__5383 (
            .O(N__30411),
            .I(measured_delay_hc_6));
    Odrv4 I__5382 (
            .O(N__30408),
            .I(measured_delay_hc_6));
    Odrv4 I__5381 (
            .O(N__30405),
            .I(measured_delay_hc_6));
    InMux I__5380 (
            .O(N__30398),
            .I(N__30395));
    LocalMux I__5379 (
            .O(N__30395),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6 ));
    CascadeMux I__5378 (
            .O(N__30392),
            .I(N__30388));
    CascadeMux I__5377 (
            .O(N__30391),
            .I(N__30384));
    InMux I__5376 (
            .O(N__30388),
            .I(N__30381));
    CascadeMux I__5375 (
            .O(N__30387),
            .I(N__30378));
    InMux I__5374 (
            .O(N__30384),
            .I(N__30375));
    LocalMux I__5373 (
            .O(N__30381),
            .I(N__30372));
    InMux I__5372 (
            .O(N__30378),
            .I(N__30369));
    LocalMux I__5371 (
            .O(N__30375),
            .I(measured_delay_hc_21));
    Odrv4 I__5370 (
            .O(N__30372),
            .I(measured_delay_hc_21));
    LocalMux I__5369 (
            .O(N__30369),
            .I(measured_delay_hc_21));
    InMux I__5368 (
            .O(N__30362),
            .I(N__30358));
    CascadeMux I__5367 (
            .O(N__30361),
            .I(N__30354));
    LocalMux I__5366 (
            .O(N__30358),
            .I(N__30350));
    InMux I__5365 (
            .O(N__30357),
            .I(N__30346));
    InMux I__5364 (
            .O(N__30354),
            .I(N__30341));
    InMux I__5363 (
            .O(N__30353),
            .I(N__30341));
    Span4Mux_v I__5362 (
            .O(N__30350),
            .I(N__30338));
    InMux I__5361 (
            .O(N__30349),
            .I(N__30335));
    LocalMux I__5360 (
            .O(N__30346),
            .I(N__30332));
    LocalMux I__5359 (
            .O(N__30341),
            .I(N__30329));
    Span4Mux_h I__5358 (
            .O(N__30338),
            .I(N__30324));
    LocalMux I__5357 (
            .O(N__30335),
            .I(N__30324));
    Span4Mux_h I__5356 (
            .O(N__30332),
            .I(N__30319));
    Span4Mux_h I__5355 (
            .O(N__30329),
            .I(N__30319));
    Odrv4 I__5354 (
            .O(N__30324),
            .I(measured_delay_hc_14));
    Odrv4 I__5353 (
            .O(N__30319),
            .I(measured_delay_hc_14));
    InMux I__5352 (
            .O(N__30314),
            .I(N__30311));
    LocalMux I__5351 (
            .O(N__30311),
            .I(N__30308));
    Odrv12 I__5350 (
            .O(N__30308),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt8 ));
    InMux I__5349 (
            .O(N__30305),
            .I(N__30302));
    LocalMux I__5348 (
            .O(N__30302),
            .I(N__30299));
    Odrv12 I__5347 (
            .O(N__30299),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    CascadeMux I__5346 (
            .O(N__30296),
            .I(N__30292));
    InMux I__5345 (
            .O(N__30295),
            .I(N__30289));
    InMux I__5344 (
            .O(N__30292),
            .I(N__30286));
    LocalMux I__5343 (
            .O(N__30289),
            .I(N__30282));
    LocalMux I__5342 (
            .O(N__30286),
            .I(N__30279));
    InMux I__5341 (
            .O(N__30285),
            .I(N__30276));
    Span4Mux_v I__5340 (
            .O(N__30282),
            .I(N__30273));
    Span4Mux_h I__5339 (
            .O(N__30279),
            .I(N__30270));
    LocalMux I__5338 (
            .O(N__30276),
            .I(N__30267));
    Span4Mux_h I__5337 (
            .O(N__30273),
            .I(N__30264));
    Span4Mux_v I__5336 (
            .O(N__30270),
            .I(N__30261));
    Odrv12 I__5335 (
            .O(N__30267),
            .I(measured_delay_hc_19));
    Odrv4 I__5334 (
            .O(N__30264),
            .I(measured_delay_hc_19));
    Odrv4 I__5333 (
            .O(N__30261),
            .I(measured_delay_hc_19));
    InMux I__5332 (
            .O(N__30254),
            .I(N__30251));
    LocalMux I__5331 (
            .O(N__30251),
            .I(N__30248));
    Span4Mux_v I__5330 (
            .O(N__30248),
            .I(N__30245));
    Odrv4 I__5329 (
            .O(N__30245),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__5328 (
            .O(N__30242),
            .I(N__30239));
    LocalMux I__5327 (
            .O(N__30239),
            .I(N__30235));
    InMux I__5326 (
            .O(N__30238),
            .I(N__30232));
    Span4Mux_h I__5325 (
            .O(N__30235),
            .I(N__30224));
    LocalMux I__5324 (
            .O(N__30232),
            .I(N__30224));
    InMux I__5323 (
            .O(N__30231),
            .I(N__30221));
    InMux I__5322 (
            .O(N__30230),
            .I(N__30218));
    InMux I__5321 (
            .O(N__30229),
            .I(N__30215));
    Span4Mux_h I__5320 (
            .O(N__30224),
            .I(N__30212));
    LocalMux I__5319 (
            .O(N__30221),
            .I(N__30209));
    LocalMux I__5318 (
            .O(N__30218),
            .I(measured_delay_hc_17));
    LocalMux I__5317 (
            .O(N__30215),
            .I(measured_delay_hc_17));
    Odrv4 I__5316 (
            .O(N__30212),
            .I(measured_delay_hc_17));
    Odrv12 I__5315 (
            .O(N__30209),
            .I(measured_delay_hc_17));
    CascadeMux I__5314 (
            .O(N__30200),
            .I(N__30197));
    InMux I__5313 (
            .O(N__30197),
            .I(N__30194));
    LocalMux I__5312 (
            .O(N__30194),
            .I(N__30191));
    Odrv12 I__5311 (
            .O(N__30191),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__5310 (
            .O(N__30188),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__5309 (
            .O(N__30185),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__5308 (
            .O(N__30182),
            .I(bfn_12_15_0_));
    InMux I__5307 (
            .O(N__30179),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__5306 (
            .O(N__30176),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__5305 (
            .O(N__30173),
            .I(N__30170));
    LocalMux I__5304 (
            .O(N__30170),
            .I(N__30167));
    Span4Mux_h I__5303 (
            .O(N__30167),
            .I(N__30164));
    Odrv4 I__5302 (
            .O(N__30164),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__5301 (
            .O(N__30161),
            .I(N__30158));
    LocalMux I__5300 (
            .O(N__30158),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__5299 (
            .O(N__30155),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ));
    CascadeMux I__5298 (
            .O(N__30152),
            .I(N__30149));
    InMux I__5297 (
            .O(N__30149),
            .I(N__30146));
    LocalMux I__5296 (
            .O(N__30146),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__5295 (
            .O(N__30143),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__5294 (
            .O(N__30140),
            .I(N__30137));
    LocalMux I__5293 (
            .O(N__30137),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__5292 (
            .O(N__30134),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ));
    CascadeMux I__5291 (
            .O(N__30131),
            .I(N__30128));
    InMux I__5290 (
            .O(N__30128),
            .I(N__30125));
    LocalMux I__5289 (
            .O(N__30125),
            .I(N__30122));
    Odrv4 I__5288 (
            .O(N__30122),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__5287 (
            .O(N__30119),
            .I(bfn_12_14_0_));
    InMux I__5286 (
            .O(N__30116),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__5285 (
            .O(N__30113),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__5284 (
            .O(N__30110),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__5283 (
            .O(N__30107),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__5282 (
            .O(N__30104),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__5281 (
            .O(N__30101),
            .I(N__30098));
    LocalMux I__5280 (
            .O(N__30098),
            .I(N__30095));
    Odrv4 I__5279 (
            .O(N__30095),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__5278 (
            .O(N__30092),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ));
    CascadeMux I__5277 (
            .O(N__30089),
            .I(N__30086));
    InMux I__5276 (
            .O(N__30086),
            .I(N__30083));
    LocalMux I__5275 (
            .O(N__30083),
            .I(N__30080));
    Odrv4 I__5274 (
            .O(N__30080),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__5273 (
            .O(N__30077),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__5272 (
            .O(N__30074),
            .I(N__30071));
    LocalMux I__5271 (
            .O(N__30071),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__5270 (
            .O(N__30068),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ));
    CascadeMux I__5269 (
            .O(N__30065),
            .I(N__30062));
    InMux I__5268 (
            .O(N__30062),
            .I(N__30059));
    LocalMux I__5267 (
            .O(N__30059),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__5266 (
            .O(N__30056),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__5265 (
            .O(N__30053),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__5264 (
            .O(N__30050),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__5263 (
            .O(N__30047),
            .I(N__30044));
    LocalMux I__5262 (
            .O(N__30044),
            .I(N__30039));
    InMux I__5261 (
            .O(N__30043),
            .I(N__30036));
    InMux I__5260 (
            .O(N__30042),
            .I(N__30033));
    Span4Mux_v I__5259 (
            .O(N__30039),
            .I(N__30028));
    LocalMux I__5258 (
            .O(N__30036),
            .I(N__30028));
    LocalMux I__5257 (
            .O(N__30033),
            .I(N__30025));
    Odrv4 I__5256 (
            .O(N__30028),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    Odrv4 I__5255 (
            .O(N__30025),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__5254 (
            .O(N__30020),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__5253 (
            .O(N__30017),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__5252 (
            .O(N__30014),
            .I(N__30010));
    InMux I__5251 (
            .O(N__30013),
            .I(N__30007));
    LocalMux I__5250 (
            .O(N__30010),
            .I(N__30001));
    LocalMux I__5249 (
            .O(N__30007),
            .I(N__30001));
    InMux I__5248 (
            .O(N__30006),
            .I(N__29998));
    Span4Mux_h I__5247 (
            .O(N__30001),
            .I(N__29995));
    LocalMux I__5246 (
            .O(N__29998),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    Odrv4 I__5245 (
            .O(N__29995),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    CascadeMux I__5244 (
            .O(N__29990),
            .I(N__29987));
    InMux I__5243 (
            .O(N__29987),
            .I(N__29984));
    LocalMux I__5242 (
            .O(N__29984),
            .I(N__29981));
    Span4Mux_h I__5241 (
            .O(N__29981),
            .I(N__29978));
    Span4Mux_h I__5240 (
            .O(N__29978),
            .I(N__29975));
    Odrv4 I__5239 (
            .O(N__29975),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__5238 (
            .O(N__29972),
            .I(N__29967));
    InMux I__5237 (
            .O(N__29971),
            .I(N__29964));
    InMux I__5236 (
            .O(N__29970),
            .I(N__29961));
    LocalMux I__5235 (
            .O(N__29967),
            .I(N__29958));
    LocalMux I__5234 (
            .O(N__29964),
            .I(N__29955));
    LocalMux I__5233 (
            .O(N__29961),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__5232 (
            .O(N__29958),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__5231 (
            .O(N__29955),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    CascadeMux I__5230 (
            .O(N__29948),
            .I(N__29945));
    InMux I__5229 (
            .O(N__29945),
            .I(N__29942));
    LocalMux I__5228 (
            .O(N__29942),
            .I(N__29939));
    Span4Mux_h I__5227 (
            .O(N__29939),
            .I(N__29936));
    Odrv4 I__5226 (
            .O(N__29936),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__5225 (
            .O(N__29933),
            .I(N__29929));
    InMux I__5224 (
            .O(N__29932),
            .I(N__29926));
    LocalMux I__5223 (
            .O(N__29929),
            .I(N__29923));
    LocalMux I__5222 (
            .O(N__29926),
            .I(N__29920));
    Odrv12 I__5221 (
            .O(N__29923),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__5220 (
            .O(N__29920),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__5219 (
            .O(N__29915),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__5218 (
            .O(N__29912),
            .I(N__29909));
    LocalMux I__5217 (
            .O(N__29909),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__5216 (
            .O(N__29906),
            .I(N__29902));
    InMux I__5215 (
            .O(N__29905),
            .I(N__29899));
    LocalMux I__5214 (
            .O(N__29902),
            .I(N__29896));
    LocalMux I__5213 (
            .O(N__29899),
            .I(N__29893));
    Odrv4 I__5212 (
            .O(N__29896),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__5211 (
            .O(N__29893),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__5210 (
            .O(N__29888),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__5209 (
            .O(N__29885),
            .I(N__29882));
    LocalMux I__5208 (
            .O(N__29882),
            .I(N__29878));
    InMux I__5207 (
            .O(N__29881),
            .I(N__29875));
    Span4Mux_v I__5206 (
            .O(N__29878),
            .I(N__29872));
    LocalMux I__5205 (
            .O(N__29875),
            .I(N__29869));
    Odrv4 I__5204 (
            .O(N__29872),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__5203 (
            .O(N__29869),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__5202 (
            .O(N__29864),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__5201 (
            .O(N__29861),
            .I(N__29857));
    InMux I__5200 (
            .O(N__29860),
            .I(N__29854));
    LocalMux I__5199 (
            .O(N__29857),
            .I(N__29851));
    LocalMux I__5198 (
            .O(N__29854),
            .I(N__29847));
    Span4Mux_h I__5197 (
            .O(N__29851),
            .I(N__29844));
    InMux I__5196 (
            .O(N__29850),
            .I(N__29841));
    Odrv12 I__5195 (
            .O(N__29847),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv4 I__5194 (
            .O(N__29844),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    LocalMux I__5193 (
            .O(N__29841),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__5192 (
            .O(N__29834),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__5191 (
            .O(N__29831),
            .I(N__29828));
    LocalMux I__5190 (
            .O(N__29828),
            .I(N__29825));
    Span4Mux_h I__5189 (
            .O(N__29825),
            .I(N__29822));
    Odrv4 I__5188 (
            .O(N__29822),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__5187 (
            .O(N__29819),
            .I(N__29815));
    InMux I__5186 (
            .O(N__29818),
            .I(N__29811));
    LocalMux I__5185 (
            .O(N__29815),
            .I(N__29808));
    InMux I__5184 (
            .O(N__29814),
            .I(N__29805));
    LocalMux I__5183 (
            .O(N__29811),
            .I(N__29802));
    Span4Mux_h I__5182 (
            .O(N__29808),
            .I(N__29799));
    LocalMux I__5181 (
            .O(N__29805),
            .I(N__29796));
    Odrv12 I__5180 (
            .O(N__29802),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__5179 (
            .O(N__29799),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__5178 (
            .O(N__29796),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__5177 (
            .O(N__29789),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__5176 (
            .O(N__29786),
            .I(N__29783));
    LocalMux I__5175 (
            .O(N__29783),
            .I(N__29780));
    Span4Mux_h I__5174 (
            .O(N__29780),
            .I(N__29777));
    Span4Mux_h I__5173 (
            .O(N__29777),
            .I(N__29774));
    Odrv4 I__5172 (
            .O(N__29774),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__5171 (
            .O(N__29771),
            .I(N__29767));
    InMux I__5170 (
            .O(N__29770),
            .I(N__29764));
    LocalMux I__5169 (
            .O(N__29767),
            .I(N__29761));
    LocalMux I__5168 (
            .O(N__29764),
            .I(N__29757));
    Span4Mux_h I__5167 (
            .O(N__29761),
            .I(N__29754));
    InMux I__5166 (
            .O(N__29760),
            .I(N__29751));
    Odrv12 I__5165 (
            .O(N__29757),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    Odrv4 I__5164 (
            .O(N__29754),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    LocalMux I__5163 (
            .O(N__29751),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__5162 (
            .O(N__29744),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__5161 (
            .O(N__29741),
            .I(N__29737));
    InMux I__5160 (
            .O(N__29740),
            .I(N__29734));
    LocalMux I__5159 (
            .O(N__29737),
            .I(N__29730));
    LocalMux I__5158 (
            .O(N__29734),
            .I(N__29727));
    InMux I__5157 (
            .O(N__29733),
            .I(N__29724));
    Span4Mux_h I__5156 (
            .O(N__29730),
            .I(N__29721));
    Span4Mux_h I__5155 (
            .O(N__29727),
            .I(N__29716));
    LocalMux I__5154 (
            .O(N__29724),
            .I(N__29716));
    Odrv4 I__5153 (
            .O(N__29721),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    Odrv4 I__5152 (
            .O(N__29716),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__5151 (
            .O(N__29711),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__5150 (
            .O(N__29708),
            .I(N__29705));
    LocalMux I__5149 (
            .O(N__29705),
            .I(N__29702));
    Span4Mux_h I__5148 (
            .O(N__29702),
            .I(N__29699));
    Odrv4 I__5147 (
            .O(N__29699),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__5146 (
            .O(N__29696),
            .I(N__29693));
    LocalMux I__5145 (
            .O(N__29693),
            .I(N__29688));
    InMux I__5144 (
            .O(N__29692),
            .I(N__29685));
    InMux I__5143 (
            .O(N__29691),
            .I(N__29682));
    Span4Mux_v I__5142 (
            .O(N__29688),
            .I(N__29675));
    LocalMux I__5141 (
            .O(N__29685),
            .I(N__29675));
    LocalMux I__5140 (
            .O(N__29682),
            .I(N__29675));
    Span4Mux_h I__5139 (
            .O(N__29675),
            .I(N__29672));
    Odrv4 I__5138 (
            .O(N__29672),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__5137 (
            .O(N__29669),
            .I(bfn_12_11_0_));
    CascadeMux I__5136 (
            .O(N__29666),
            .I(N__29663));
    InMux I__5135 (
            .O(N__29663),
            .I(N__29660));
    LocalMux I__5134 (
            .O(N__29660),
            .I(N__29657));
    Span4Mux_v I__5133 (
            .O(N__29657),
            .I(N__29654));
    Odrv4 I__5132 (
            .O(N__29654),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    InMux I__5131 (
            .O(N__29651),
            .I(N__29647));
    InMux I__5130 (
            .O(N__29650),
            .I(N__29643));
    LocalMux I__5129 (
            .O(N__29647),
            .I(N__29640));
    InMux I__5128 (
            .O(N__29646),
            .I(N__29637));
    LocalMux I__5127 (
            .O(N__29643),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    Odrv4 I__5126 (
            .O(N__29640),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    LocalMux I__5125 (
            .O(N__29637),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    InMux I__5124 (
            .O(N__29630),
            .I(N__29626));
    InMux I__5123 (
            .O(N__29629),
            .I(N__29622));
    LocalMux I__5122 (
            .O(N__29626),
            .I(N__29619));
    InMux I__5121 (
            .O(N__29625),
            .I(N__29616));
    LocalMux I__5120 (
            .O(N__29622),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    Odrv4 I__5119 (
            .O(N__29619),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    LocalMux I__5118 (
            .O(N__29616),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    InMux I__5117 (
            .O(N__29609),
            .I(N__29605));
    InMux I__5116 (
            .O(N__29608),
            .I(N__29601));
    LocalMux I__5115 (
            .O(N__29605),
            .I(N__29598));
    InMux I__5114 (
            .O(N__29604),
            .I(N__29595));
    LocalMux I__5113 (
            .O(N__29601),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    Odrv4 I__5112 (
            .O(N__29598),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    LocalMux I__5111 (
            .O(N__29595),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__5110 (
            .O(N__29588),
            .I(N__29585));
    LocalMux I__5109 (
            .O(N__29585),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__5108 (
            .O(N__29582),
            .I(N__29579));
    LocalMux I__5107 (
            .O(N__29579),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__5106 (
            .O(N__29576),
            .I(N__29573));
    LocalMux I__5105 (
            .O(N__29573),
            .I(N__29570));
    Span4Mux_v I__5104 (
            .O(N__29570),
            .I(N__29565));
    InMux I__5103 (
            .O(N__29569),
            .I(N__29562));
    InMux I__5102 (
            .O(N__29568),
            .I(N__29559));
    Span4Mux_v I__5101 (
            .O(N__29565),
            .I(N__29556));
    LocalMux I__5100 (
            .O(N__29562),
            .I(N__29553));
    LocalMux I__5099 (
            .O(N__29559),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv4 I__5098 (
            .O(N__29556),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv12 I__5097 (
            .O(N__29553),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    InMux I__5096 (
            .O(N__29546),
            .I(N__29543));
    LocalMux I__5095 (
            .O(N__29543),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    InMux I__5094 (
            .O(N__29540),
            .I(N__29537));
    LocalMux I__5093 (
            .O(N__29537),
            .I(N__29534));
    Span4Mux_h I__5092 (
            .O(N__29534),
            .I(N__29531));
    Odrv4 I__5091 (
            .O(N__29531),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ));
    InMux I__5090 (
            .O(N__29528),
            .I(N__29525));
    LocalMux I__5089 (
            .O(N__29525),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    CascadeMux I__5088 (
            .O(N__29522),
            .I(N__29519));
    InMux I__5087 (
            .O(N__29519),
            .I(N__29513));
    InMux I__5086 (
            .O(N__29518),
            .I(N__29510));
    CascadeMux I__5085 (
            .O(N__29517),
            .I(N__29507));
    InMux I__5084 (
            .O(N__29516),
            .I(N__29504));
    LocalMux I__5083 (
            .O(N__29513),
            .I(N__29498));
    LocalMux I__5082 (
            .O(N__29510),
            .I(N__29498));
    InMux I__5081 (
            .O(N__29507),
            .I(N__29495));
    LocalMux I__5080 (
            .O(N__29504),
            .I(N__29492));
    CascadeMux I__5079 (
            .O(N__29503),
            .I(N__29489));
    Span4Mux_h I__5078 (
            .O(N__29498),
            .I(N__29486));
    LocalMux I__5077 (
            .O(N__29495),
            .I(N__29483));
    Span4Mux_h I__5076 (
            .O(N__29492),
            .I(N__29480));
    InMux I__5075 (
            .O(N__29489),
            .I(N__29477));
    Span4Mux_v I__5074 (
            .O(N__29486),
            .I(N__29474));
    Odrv4 I__5073 (
            .O(N__29483),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__5072 (
            .O(N__29480),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__5071 (
            .O(N__29477),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__5070 (
            .O(N__29474),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__5069 (
            .O(N__29465),
            .I(N__29462));
    InMux I__5068 (
            .O(N__29462),
            .I(N__29459));
    LocalMux I__5067 (
            .O(N__29459),
            .I(N__29456));
    Span4Mux_v I__5066 (
            .O(N__29456),
            .I(N__29453));
    Span4Mux_v I__5065 (
            .O(N__29453),
            .I(N__29450));
    Odrv4 I__5064 (
            .O(N__29450),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    CascadeMux I__5063 (
            .O(N__29447),
            .I(N__29444));
    InMux I__5062 (
            .O(N__29444),
            .I(N__29441));
    LocalMux I__5061 (
            .O(N__29441),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__5060 (
            .O(N__29438),
            .I(N__29435));
    LocalMux I__5059 (
            .O(N__29435),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    InMux I__5058 (
            .O(N__29432),
            .I(N__29429));
    LocalMux I__5057 (
            .O(N__29429),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__5056 (
            .O(N__29426),
            .I(N__29423));
    LocalMux I__5055 (
            .O(N__29423),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    InMux I__5054 (
            .O(N__29420),
            .I(N__29417));
    LocalMux I__5053 (
            .O(N__29417),
            .I(\delay_measurement_inst.N_59 ));
    InMux I__5052 (
            .O(N__29414),
            .I(N__29406));
    InMux I__5051 (
            .O(N__29413),
            .I(N__29395));
    InMux I__5050 (
            .O(N__29412),
            .I(N__29395));
    InMux I__5049 (
            .O(N__29411),
            .I(N__29395));
    InMux I__5048 (
            .O(N__29410),
            .I(N__29395));
    InMux I__5047 (
            .O(N__29409),
            .I(N__29395));
    LocalMux I__5046 (
            .O(N__29406),
            .I(\delay_measurement_inst.N_270 ));
    LocalMux I__5045 (
            .O(N__29395),
            .I(\delay_measurement_inst.N_270 ));
    CascadeMux I__5044 (
            .O(N__29390),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_ ));
    CascadeMux I__5043 (
            .O(N__29387),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7_cascade_ ));
    InMux I__5042 (
            .O(N__29384),
            .I(N__29381));
    LocalMux I__5041 (
            .O(N__29381),
            .I(N__29378));
    Span4Mux_h I__5040 (
            .O(N__29378),
            .I(N__29375));
    Odrv4 I__5039 (
            .O(N__29375),
            .I(delay_tr_input_c));
    InMux I__5038 (
            .O(N__29372),
            .I(N__29369));
    LocalMux I__5037 (
            .O(N__29369),
            .I(delay_tr_d1));
    InMux I__5036 (
            .O(N__29366),
            .I(N__29360));
    InMux I__5035 (
            .O(N__29365),
            .I(N__29355));
    InMux I__5034 (
            .O(N__29364),
            .I(N__29355));
    InMux I__5033 (
            .O(N__29363),
            .I(N__29352));
    LocalMux I__5032 (
            .O(N__29360),
            .I(delay_tr_d2));
    LocalMux I__5031 (
            .O(N__29355),
            .I(delay_tr_d2));
    LocalMux I__5030 (
            .O(N__29352),
            .I(delay_tr_d2));
    InMux I__5029 (
            .O(N__29345),
            .I(N__29340));
    InMux I__5028 (
            .O(N__29344),
            .I(N__29337));
    InMux I__5027 (
            .O(N__29343),
            .I(N__29334));
    LocalMux I__5026 (
            .O(N__29340),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__5025 (
            .O(N__29337),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__5024 (
            .O(N__29334),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__5023 (
            .O(N__29327),
            .I(N__29322));
    InMux I__5022 (
            .O(N__29326),
            .I(N__29319));
    InMux I__5021 (
            .O(N__29325),
            .I(N__29316));
    LocalMux I__5020 (
            .O(N__29322),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__5019 (
            .O(N__29319),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__5018 (
            .O(N__29316),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__5017 (
            .O(N__29309),
            .I(N__29306));
    LocalMux I__5016 (
            .O(N__29306),
            .I(N__29302));
    InMux I__5015 (
            .O(N__29305),
            .I(N__29299));
    Span4Mux_v I__5014 (
            .O(N__29302),
            .I(N__29294));
    LocalMux I__5013 (
            .O(N__29299),
            .I(N__29294));
    Span4Mux_v I__5012 (
            .O(N__29294),
            .I(N__29291));
    Span4Mux_v I__5011 (
            .O(N__29291),
            .I(N__29288));
    Span4Mux_v I__5010 (
            .O(N__29288),
            .I(N__29285));
    Odrv4 I__5009 (
            .O(N__29285),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__5008 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__5007 (
            .O(N__29279),
            .I(N__29275));
    InMux I__5006 (
            .O(N__29278),
            .I(N__29272));
    Span4Mux_v I__5005 (
            .O(N__29275),
            .I(N__29268));
    LocalMux I__5004 (
            .O(N__29272),
            .I(N__29265));
    InMux I__5003 (
            .O(N__29271),
            .I(N__29262));
    Span4Mux_v I__5002 (
            .O(N__29268),
            .I(N__29259));
    Span4Mux_h I__5001 (
            .O(N__29265),
            .I(N__29256));
    LocalMux I__5000 (
            .O(N__29262),
            .I(N__29253));
    Sp12to4 I__4999 (
            .O(N__29259),
            .I(N__29250));
    Sp12to4 I__4998 (
            .O(N__29256),
            .I(N__29245));
    Sp12to4 I__4997 (
            .O(N__29253),
            .I(N__29245));
    Span12Mux_h I__4996 (
            .O(N__29250),
            .I(N__29240));
    Span12Mux_v I__4995 (
            .O(N__29245),
            .I(N__29240));
    Odrv12 I__4994 (
            .O(N__29240),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__4993 (
            .O(N__29237),
            .I(N__29231));
    InMux I__4992 (
            .O(N__29236),
            .I(N__29231));
    LocalMux I__4991 (
            .O(N__29231),
            .I(N__29228));
    Span4Mux_v I__4990 (
            .O(N__29228),
            .I(N__29223));
    InMux I__4989 (
            .O(N__29227),
            .I(N__29220));
    InMux I__4988 (
            .O(N__29226),
            .I(N__29217));
    Span4Mux_h I__4987 (
            .O(N__29223),
            .I(N__29214));
    LocalMux I__4986 (
            .O(N__29220),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4985 (
            .O(N__29217),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__4984 (
            .O(N__29214),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    CascadeMux I__4983 (
            .O(N__29207),
            .I(N__29204));
    InMux I__4982 (
            .O(N__29204),
            .I(N__29200));
    InMux I__4981 (
            .O(N__29203),
            .I(N__29197));
    LocalMux I__4980 (
            .O(N__29200),
            .I(N__29192));
    LocalMux I__4979 (
            .O(N__29197),
            .I(N__29192));
    Odrv12 I__4978 (
            .O(N__29192),
            .I(measured_delay_hc_25));
    CascadeMux I__4977 (
            .O(N__29189),
            .I(N__29186));
    InMux I__4976 (
            .O(N__29186),
            .I(N__29182));
    InMux I__4975 (
            .O(N__29185),
            .I(N__29179));
    LocalMux I__4974 (
            .O(N__29182),
            .I(measured_delay_hc_24));
    LocalMux I__4973 (
            .O(N__29179),
            .I(measured_delay_hc_24));
    CascadeMux I__4972 (
            .O(N__29174),
            .I(N__29171));
    InMux I__4971 (
            .O(N__29171),
            .I(N__29167));
    InMux I__4970 (
            .O(N__29170),
            .I(N__29164));
    LocalMux I__4969 (
            .O(N__29167),
            .I(N__29161));
    LocalMux I__4968 (
            .O(N__29164),
            .I(measured_delay_hc_26));
    Odrv4 I__4967 (
            .O(N__29161),
            .I(measured_delay_hc_26));
    CascadeMux I__4966 (
            .O(N__29156),
            .I(N__29153));
    InMux I__4965 (
            .O(N__29153),
            .I(N__29149));
    InMux I__4964 (
            .O(N__29152),
            .I(N__29146));
    LocalMux I__4963 (
            .O(N__29149),
            .I(measured_delay_hc_23));
    LocalMux I__4962 (
            .O(N__29146),
            .I(measured_delay_hc_23));
    InMux I__4961 (
            .O(N__29141),
            .I(N__29138));
    LocalMux I__4960 (
            .O(N__29138),
            .I(N__29134));
    InMux I__4959 (
            .O(N__29137),
            .I(N__29131));
    Span4Mux_h I__4958 (
            .O(N__29134),
            .I(N__29128));
    LocalMux I__4957 (
            .O(N__29131),
            .I(measured_delay_hc_28));
    Odrv4 I__4956 (
            .O(N__29128),
            .I(measured_delay_hc_28));
    CascadeMux I__4955 (
            .O(N__29123),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4_cascade_ ));
    InMux I__4954 (
            .O(N__29120),
            .I(N__29116));
    CascadeMux I__4953 (
            .O(N__29119),
            .I(N__29113));
    LocalMux I__4952 (
            .O(N__29116),
            .I(N__29110));
    InMux I__4951 (
            .O(N__29113),
            .I(N__29107));
    Odrv4 I__4950 (
            .O(N__29110),
            .I(\delay_measurement_inst.elapsed_time_hc_30 ));
    LocalMux I__4949 (
            .O(N__29107),
            .I(\delay_measurement_inst.elapsed_time_hc_30 ));
    InMux I__4948 (
            .O(N__29102),
            .I(N__29099));
    LocalMux I__4947 (
            .O(N__29099),
            .I(\delay_measurement_inst.N_51 ));
    InMux I__4946 (
            .O(N__29096),
            .I(N__29093));
    LocalMux I__4945 (
            .O(N__29093),
            .I(N__29089));
    InMux I__4944 (
            .O(N__29092),
            .I(N__29086));
    Odrv4 I__4943 (
            .O(N__29089),
            .I(measured_delay_hc_27));
    LocalMux I__4942 (
            .O(N__29086),
            .I(measured_delay_hc_27));
    InMux I__4941 (
            .O(N__29081),
            .I(N__29078));
    LocalMux I__4940 (
            .O(N__29078),
            .I(\delay_measurement_inst.N_25 ));
    IoInMux I__4939 (
            .O(N__29075),
            .I(N__29072));
    LocalMux I__4938 (
            .O(N__29072),
            .I(\delay_measurement_inst.delay_tr_timer.N_304_i ));
    CascadeMux I__4937 (
            .O(N__29069),
            .I(\delay_measurement_inst.N_33_cascade_ ));
    InMux I__4936 (
            .O(N__29066),
            .I(N__29063));
    LocalMux I__4935 (
            .O(N__29063),
            .I(N__29060));
    Odrv12 I__4934 (
            .O(N__29060),
            .I(\delay_measurement_inst.N_38 ));
    InMux I__4933 (
            .O(N__29057),
            .I(N__29054));
    LocalMux I__4932 (
            .O(N__29054),
            .I(N__29049));
    InMux I__4931 (
            .O(N__29053),
            .I(N__29044));
    InMux I__4930 (
            .O(N__29052),
            .I(N__29044));
    Odrv12 I__4929 (
            .O(N__29049),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__4928 (
            .O(N__29044),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    InMux I__4927 (
            .O(N__29039),
            .I(N__29036));
    LocalMux I__4926 (
            .O(N__29036),
            .I(N__29032));
    InMux I__4925 (
            .O(N__29035),
            .I(N__29029));
    Span4Mux_v I__4924 (
            .O(N__29032),
            .I(N__29026));
    LocalMux I__4923 (
            .O(N__29029),
            .I(N__29023));
    Odrv4 I__4922 (
            .O(N__29026),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__4921 (
            .O(N__29023),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__4920 (
            .O(N__29018),
            .I(N__29014));
    InMux I__4919 (
            .O(N__29017),
            .I(N__29011));
    LocalMux I__4918 (
            .O(N__29014),
            .I(N__29008));
    LocalMux I__4917 (
            .O(N__29011),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ));
    Odrv4 I__4916 (
            .O(N__29008),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ));
    CascadeMux I__4915 (
            .O(N__29003),
            .I(N__29000));
    InMux I__4914 (
            .O(N__29000),
            .I(N__28997));
    LocalMux I__4913 (
            .O(N__28997),
            .I(N__28994));
    Odrv4 I__4912 (
            .O(N__28994),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_0 ));
    InMux I__4911 (
            .O(N__28991),
            .I(N__28988));
    LocalMux I__4910 (
            .O(N__28988),
            .I(N__28985));
    Odrv4 I__4909 (
            .O(N__28985),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ));
    InMux I__4908 (
            .O(N__28982),
            .I(N__28978));
    InMux I__4907 (
            .O(N__28981),
            .I(N__28974));
    LocalMux I__4906 (
            .O(N__28978),
            .I(N__28971));
    CascadeMux I__4905 (
            .O(N__28977),
            .I(N__28968));
    LocalMux I__4904 (
            .O(N__28974),
            .I(N__28965));
    Span4Mux_h I__4903 (
            .O(N__28971),
            .I(N__28962));
    InMux I__4902 (
            .O(N__28968),
            .I(N__28959));
    Span4Mux_h I__4901 (
            .O(N__28965),
            .I(N__28956));
    Odrv4 I__4900 (
            .O(N__28962),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__4899 (
            .O(N__28959),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    Odrv4 I__4898 (
            .O(N__28956),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    CEMux I__4897 (
            .O(N__28949),
            .I(N__28945));
    CEMux I__4896 (
            .O(N__28948),
            .I(N__28941));
    LocalMux I__4895 (
            .O(N__28945),
            .I(N__28937));
    CEMux I__4894 (
            .O(N__28944),
            .I(N__28934));
    LocalMux I__4893 (
            .O(N__28941),
            .I(N__28931));
    CEMux I__4892 (
            .O(N__28940),
            .I(N__28928));
    Span4Mux_v I__4891 (
            .O(N__28937),
            .I(N__28923));
    LocalMux I__4890 (
            .O(N__28934),
            .I(N__28923));
    Span4Mux_v I__4889 (
            .O(N__28931),
            .I(N__28918));
    LocalMux I__4888 (
            .O(N__28928),
            .I(N__28918));
    Sp12to4 I__4887 (
            .O(N__28923),
            .I(N__28915));
    Odrv4 I__4886 (
            .O(N__28918),
            .I(\delay_measurement_inst.delay_hc_timer.N_303_i ));
    Odrv12 I__4885 (
            .O(N__28915),
            .I(\delay_measurement_inst.delay_hc_timer.N_303_i ));
    InMux I__4884 (
            .O(N__28910),
            .I(N__28907));
    LocalMux I__4883 (
            .O(N__28907),
            .I(N__28904));
    Odrv4 I__4882 (
            .O(N__28904),
            .I(\delay_measurement_inst.N_28 ));
    InMux I__4881 (
            .O(N__28901),
            .I(N__28896));
    InMux I__4880 (
            .O(N__28900),
            .I(N__28893));
    InMux I__4879 (
            .O(N__28899),
            .I(N__28890));
    LocalMux I__4878 (
            .O(N__28896),
            .I(N__28885));
    LocalMux I__4877 (
            .O(N__28893),
            .I(N__28885));
    LocalMux I__4876 (
            .O(N__28890),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv12 I__4875 (
            .O(N__28885),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__4874 (
            .O(N__28880),
            .I(N__28877));
    LocalMux I__4873 (
            .O(N__28877),
            .I(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ));
    CascadeMux I__4872 (
            .O(N__28874),
            .I(N__28871));
    InMux I__4871 (
            .O(N__28871),
            .I(N__28868));
    LocalMux I__4870 (
            .O(N__28868),
            .I(N__28865));
    Span4Mux_h I__4869 (
            .O(N__28865),
            .I(N__28862));
    Odrv4 I__4868 (
            .O(N__28862),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__4867 (
            .O(N__28859),
            .I(N__28856));
    InMux I__4866 (
            .O(N__28856),
            .I(N__28853));
    LocalMux I__4865 (
            .O(N__28853),
            .I(N__28850));
    Odrv12 I__4864 (
            .O(N__28850),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CEMux I__4863 (
            .O(N__28847),
            .I(N__28844));
    LocalMux I__4862 (
            .O(N__28844),
            .I(N__28839));
    CEMux I__4861 (
            .O(N__28843),
            .I(N__28836));
    CEMux I__4860 (
            .O(N__28842),
            .I(N__28833));
    Span4Mux_h I__4859 (
            .O(N__28839),
            .I(N__28828));
    LocalMux I__4858 (
            .O(N__28836),
            .I(N__28825));
    LocalMux I__4857 (
            .O(N__28833),
            .I(N__28822));
    CEMux I__4856 (
            .O(N__28832),
            .I(N__28819));
    CEMux I__4855 (
            .O(N__28831),
            .I(N__28816));
    Span4Mux_v I__4854 (
            .O(N__28828),
            .I(N__28813));
    Span4Mux_h I__4853 (
            .O(N__28825),
            .I(N__28810));
    Span4Mux_v I__4852 (
            .O(N__28822),
            .I(N__28807));
    LocalMux I__4851 (
            .O(N__28819),
            .I(N__28802));
    LocalMux I__4850 (
            .O(N__28816),
            .I(N__28802));
    Odrv4 I__4849 (
            .O(N__28813),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__4848 (
            .O(N__28810),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__4847 (
            .O(N__28807),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv12 I__4846 (
            .O(N__28802),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__4845 (
            .O(N__28793),
            .I(N__28790));
    LocalMux I__4844 (
            .O(N__28790),
            .I(N__28786));
    CascadeMux I__4843 (
            .O(N__28789),
            .I(N__28783));
    Span4Mux_h I__4842 (
            .O(N__28786),
            .I(N__28780));
    InMux I__4841 (
            .O(N__28783),
            .I(N__28777));
    Span4Mux_v I__4840 (
            .O(N__28780),
            .I(N__28774));
    LocalMux I__4839 (
            .O(N__28777),
            .I(N__28771));
    Span4Mux_v I__4838 (
            .O(N__28774),
            .I(N__28768));
    Odrv4 I__4837 (
            .O(N__28771),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    Odrv4 I__4836 (
            .O(N__28768),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__4835 (
            .O(N__28763),
            .I(N__28760));
    LocalMux I__4834 (
            .O(N__28760),
            .I(N__28754));
    InMux I__4833 (
            .O(N__28759),
            .I(N__28747));
    InMux I__4832 (
            .O(N__28758),
            .I(N__28747));
    InMux I__4831 (
            .O(N__28757),
            .I(N__28747));
    Odrv4 I__4830 (
            .O(N__28754),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__4829 (
            .O(N__28747),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__4828 (
            .O(N__28742),
            .I(N__28739));
    LocalMux I__4827 (
            .O(N__28739),
            .I(N__28736));
    Odrv4 I__4826 (
            .O(N__28736),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    CascadeMux I__4825 (
            .O(N__28733),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ));
    InMux I__4824 (
            .O(N__28730),
            .I(N__28726));
    InMux I__4823 (
            .O(N__28729),
            .I(N__28722));
    LocalMux I__4822 (
            .O(N__28726),
            .I(N__28719));
    InMux I__4821 (
            .O(N__28725),
            .I(N__28716));
    LocalMux I__4820 (
            .O(N__28722),
            .I(N__28713));
    Span4Mux_v I__4819 (
            .O(N__28719),
            .I(N__28708));
    LocalMux I__4818 (
            .O(N__28716),
            .I(N__28705));
    Span4Mux_h I__4817 (
            .O(N__28713),
            .I(N__28702));
    InMux I__4816 (
            .O(N__28712),
            .I(N__28697));
    InMux I__4815 (
            .O(N__28711),
            .I(N__28697));
    Odrv4 I__4814 (
            .O(N__28708),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__4813 (
            .O(N__28705),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__4812 (
            .O(N__28702),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__4811 (
            .O(N__28697),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__4810 (
            .O(N__28688),
            .I(N__28685));
    LocalMux I__4809 (
            .O(N__28685),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ));
    CascadeMux I__4808 (
            .O(N__28682),
            .I(N__28678));
    CascadeMux I__4807 (
            .O(N__28681),
            .I(N__28674));
    InMux I__4806 (
            .O(N__28678),
            .I(N__28667));
    InMux I__4805 (
            .O(N__28677),
            .I(N__28667));
    InMux I__4804 (
            .O(N__28674),
            .I(N__28667));
    LocalMux I__4803 (
            .O(N__28667),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_16 ));
    CascadeMux I__4802 (
            .O(N__28664),
            .I(N__28655));
    CascadeMux I__4801 (
            .O(N__28663),
            .I(N__28651));
    CascadeMux I__4800 (
            .O(N__28662),
            .I(N__28647));
    CascadeMux I__4799 (
            .O(N__28661),
            .I(N__28643));
    CascadeMux I__4798 (
            .O(N__28660),
            .I(N__28639));
    CascadeMux I__4797 (
            .O(N__28659),
            .I(N__28635));
    InMux I__4796 (
            .O(N__28658),
            .I(N__28624));
    InMux I__4795 (
            .O(N__28655),
            .I(N__28624));
    InMux I__4794 (
            .O(N__28654),
            .I(N__28624));
    InMux I__4793 (
            .O(N__28651),
            .I(N__28624));
    InMux I__4792 (
            .O(N__28650),
            .I(N__28607));
    InMux I__4791 (
            .O(N__28647),
            .I(N__28607));
    InMux I__4790 (
            .O(N__28646),
            .I(N__28607));
    InMux I__4789 (
            .O(N__28643),
            .I(N__28607));
    InMux I__4788 (
            .O(N__28642),
            .I(N__28607));
    InMux I__4787 (
            .O(N__28639),
            .I(N__28607));
    InMux I__4786 (
            .O(N__28638),
            .I(N__28607));
    InMux I__4785 (
            .O(N__28635),
            .I(N__28607));
    CascadeMux I__4784 (
            .O(N__28634),
            .I(N__28603));
    CascadeMux I__4783 (
            .O(N__28633),
            .I(N__28599));
    LocalMux I__4782 (
            .O(N__28624),
            .I(N__28594));
    LocalMux I__4781 (
            .O(N__28607),
            .I(N__28594));
    InMux I__4780 (
            .O(N__28606),
            .I(N__28585));
    InMux I__4779 (
            .O(N__28603),
            .I(N__28585));
    InMux I__4778 (
            .O(N__28602),
            .I(N__28585));
    InMux I__4777 (
            .O(N__28599),
            .I(N__28585));
    Span4Mux_v I__4776 (
            .O(N__28594),
            .I(N__28580));
    LocalMux I__4775 (
            .O(N__28585),
            .I(N__28580));
    Span4Mux_h I__4774 (
            .O(N__28580),
            .I(N__28577));
    Odrv4 I__4773 (
            .O(N__28577),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__4772 (
            .O(N__28574),
            .I(N__28570));
    InMux I__4771 (
            .O(N__28573),
            .I(N__28566));
    LocalMux I__4770 (
            .O(N__28570),
            .I(N__28563));
    InMux I__4769 (
            .O(N__28569),
            .I(N__28560));
    LocalMux I__4768 (
            .O(N__28566),
            .I(N__28557));
    Span4Mux_v I__4767 (
            .O(N__28563),
            .I(N__28554));
    LocalMux I__4766 (
            .O(N__28560),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__4765 (
            .O(N__28557),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__4764 (
            .O(N__28554),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__4763 (
            .O(N__28547),
            .I(N__28542));
    InMux I__4762 (
            .O(N__28546),
            .I(N__28539));
    InMux I__4761 (
            .O(N__28545),
            .I(N__28536));
    LocalMux I__4760 (
            .O(N__28542),
            .I(N__28533));
    LocalMux I__4759 (
            .O(N__28539),
            .I(N__28530));
    LocalMux I__4758 (
            .O(N__28536),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__4757 (
            .O(N__28533),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv12 I__4756 (
            .O(N__28530),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    InMux I__4755 (
            .O(N__28523),
            .I(N__28519));
    InMux I__4754 (
            .O(N__28522),
            .I(N__28516));
    LocalMux I__4753 (
            .O(N__28519),
            .I(N__28510));
    LocalMux I__4752 (
            .O(N__28516),
            .I(N__28510));
    InMux I__4751 (
            .O(N__28515),
            .I(N__28507));
    Span4Mux_v I__4750 (
            .O(N__28510),
            .I(N__28504));
    LocalMux I__4749 (
            .O(N__28507),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    Odrv4 I__4748 (
            .O(N__28504),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    CascadeMux I__4747 (
            .O(N__28499),
            .I(N__28495));
    InMux I__4746 (
            .O(N__28498),
            .I(N__28492));
    InMux I__4745 (
            .O(N__28495),
            .I(N__28488));
    LocalMux I__4744 (
            .O(N__28492),
            .I(N__28485));
    InMux I__4743 (
            .O(N__28491),
            .I(N__28482));
    LocalMux I__4742 (
            .O(N__28488),
            .I(N__28477));
    Span4Mux_h I__4741 (
            .O(N__28485),
            .I(N__28477));
    LocalMux I__4740 (
            .O(N__28482),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    Odrv4 I__4739 (
            .O(N__28477),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    CascadeMux I__4738 (
            .O(N__28472),
            .I(N__28468));
    InMux I__4737 (
            .O(N__28471),
            .I(N__28465));
    InMux I__4736 (
            .O(N__28468),
            .I(N__28460));
    LocalMux I__4735 (
            .O(N__28465),
            .I(N__28457));
    InMux I__4734 (
            .O(N__28464),
            .I(N__28454));
    InMux I__4733 (
            .O(N__28463),
            .I(N__28451));
    LocalMux I__4732 (
            .O(N__28460),
            .I(N__28447));
    Span4Mux_v I__4731 (
            .O(N__28457),
            .I(N__28442));
    LocalMux I__4730 (
            .O(N__28454),
            .I(N__28442));
    LocalMux I__4729 (
            .O(N__28451),
            .I(N__28439));
    InMux I__4728 (
            .O(N__28450),
            .I(N__28436));
    Span4Mux_v I__4727 (
            .O(N__28447),
            .I(N__28431));
    Span4Mux_h I__4726 (
            .O(N__28442),
            .I(N__28431));
    Odrv4 I__4725 (
            .O(N__28439),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__4724 (
            .O(N__28436),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__4723 (
            .O(N__28431),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__4722 (
            .O(N__28424),
            .I(N__28421));
    LocalMux I__4721 (
            .O(N__28421),
            .I(N__28418));
    Span4Mux_v I__4720 (
            .O(N__28418),
            .I(N__28415));
    Odrv4 I__4719 (
            .O(N__28415),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    InMux I__4718 (
            .O(N__28412),
            .I(N__28409));
    LocalMux I__4717 (
            .O(N__28409),
            .I(N__28406));
    Odrv4 I__4716 (
            .O(N__28406),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ));
    InMux I__4715 (
            .O(N__28403),
            .I(N__28400));
    LocalMux I__4714 (
            .O(N__28400),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__4713 (
            .O(N__28397),
            .I(N__28393));
    InMux I__4712 (
            .O(N__28396),
            .I(N__28389));
    LocalMux I__4711 (
            .O(N__28393),
            .I(N__28386));
    InMux I__4710 (
            .O(N__28392),
            .I(N__28383));
    LocalMux I__4709 (
            .O(N__28389),
            .I(N__28380));
    Span4Mux_v I__4708 (
            .O(N__28386),
            .I(N__28375));
    LocalMux I__4707 (
            .O(N__28383),
            .I(N__28375));
    Span4Mux_h I__4706 (
            .O(N__28380),
            .I(N__28371));
    Span4Mux_h I__4705 (
            .O(N__28375),
            .I(N__28368));
    InMux I__4704 (
            .O(N__28374),
            .I(N__28365));
    Odrv4 I__4703 (
            .O(N__28371),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__4702 (
            .O(N__28368),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__4701 (
            .O(N__28365),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__4700 (
            .O(N__28358),
            .I(N__28355));
    LocalMux I__4699 (
            .O(N__28355),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    CascadeMux I__4698 (
            .O(N__28352),
            .I(N__28348));
    CascadeMux I__4697 (
            .O(N__28351),
            .I(N__28344));
    InMux I__4696 (
            .O(N__28348),
            .I(N__28341));
    InMux I__4695 (
            .O(N__28347),
            .I(N__28338));
    InMux I__4694 (
            .O(N__28344),
            .I(N__28335));
    LocalMux I__4693 (
            .O(N__28341),
            .I(N__28332));
    LocalMux I__4692 (
            .O(N__28338),
            .I(N__28327));
    LocalMux I__4691 (
            .O(N__28335),
            .I(N__28327));
    Span4Mux_v I__4690 (
            .O(N__28332),
            .I(N__28323));
    Span4Mux_v I__4689 (
            .O(N__28327),
            .I(N__28320));
    InMux I__4688 (
            .O(N__28326),
            .I(N__28317));
    Odrv4 I__4687 (
            .O(N__28323),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4686 (
            .O(N__28320),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__4685 (
            .O(N__28317),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__4684 (
            .O(N__28310),
            .I(N__28307));
    LocalMux I__4683 (
            .O(N__28307),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__4682 (
            .O(N__28304),
            .I(N__28289));
    CascadeMux I__4681 (
            .O(N__28303),
            .I(N__28286));
    InMux I__4680 (
            .O(N__28302),
            .I(N__28274));
    InMux I__4679 (
            .O(N__28301),
            .I(N__28274));
    InMux I__4678 (
            .O(N__28300),
            .I(N__28269));
    InMux I__4677 (
            .O(N__28299),
            .I(N__28269));
    InMux I__4676 (
            .O(N__28298),
            .I(N__28266));
    InMux I__4675 (
            .O(N__28297),
            .I(N__28255));
    InMux I__4674 (
            .O(N__28296),
            .I(N__28255));
    InMux I__4673 (
            .O(N__28295),
            .I(N__28255));
    InMux I__4672 (
            .O(N__28294),
            .I(N__28255));
    InMux I__4671 (
            .O(N__28293),
            .I(N__28255));
    CascadeMux I__4670 (
            .O(N__28292),
            .I(N__28243));
    InMux I__4669 (
            .O(N__28289),
            .I(N__28230));
    InMux I__4668 (
            .O(N__28286),
            .I(N__28230));
    InMux I__4667 (
            .O(N__28285),
            .I(N__28230));
    InMux I__4666 (
            .O(N__28284),
            .I(N__28230));
    InMux I__4665 (
            .O(N__28283),
            .I(N__28230));
    InMux I__4664 (
            .O(N__28282),
            .I(N__28221));
    InMux I__4663 (
            .O(N__28281),
            .I(N__28221));
    InMux I__4662 (
            .O(N__28280),
            .I(N__28221));
    InMux I__4661 (
            .O(N__28279),
            .I(N__28221));
    LocalMux I__4660 (
            .O(N__28274),
            .I(N__28216));
    LocalMux I__4659 (
            .O(N__28269),
            .I(N__28216));
    LocalMux I__4658 (
            .O(N__28266),
            .I(N__28213));
    LocalMux I__4657 (
            .O(N__28255),
            .I(N__28210));
    InMux I__4656 (
            .O(N__28254),
            .I(N__28205));
    InMux I__4655 (
            .O(N__28253),
            .I(N__28205));
    InMux I__4654 (
            .O(N__28252),
            .I(N__28196));
    InMux I__4653 (
            .O(N__28251),
            .I(N__28196));
    InMux I__4652 (
            .O(N__28250),
            .I(N__28196));
    InMux I__4651 (
            .O(N__28249),
            .I(N__28196));
    InMux I__4650 (
            .O(N__28248),
            .I(N__28183));
    InMux I__4649 (
            .O(N__28247),
            .I(N__28183));
    InMux I__4648 (
            .O(N__28246),
            .I(N__28183));
    InMux I__4647 (
            .O(N__28243),
            .I(N__28183));
    InMux I__4646 (
            .O(N__28242),
            .I(N__28183));
    InMux I__4645 (
            .O(N__28241),
            .I(N__28183));
    LocalMux I__4644 (
            .O(N__28230),
            .I(N__28178));
    LocalMux I__4643 (
            .O(N__28221),
            .I(N__28178));
    Span4Mux_h I__4642 (
            .O(N__28216),
            .I(N__28173));
    Span4Mux_h I__4641 (
            .O(N__28213),
            .I(N__28173));
    Span4Mux_v I__4640 (
            .O(N__28210),
            .I(N__28170));
    LocalMux I__4639 (
            .O(N__28205),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__4638 (
            .O(N__28196),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__4637 (
            .O(N__28183),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__4636 (
            .O(N__28178),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__4635 (
            .O(N__28173),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__4634 (
            .O(N__28170),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__4633 (
            .O(N__28157),
            .I(N__28133));
    InMux I__4632 (
            .O(N__28156),
            .I(N__28133));
    InMux I__4631 (
            .O(N__28155),
            .I(N__28133));
    InMux I__4630 (
            .O(N__28154),
            .I(N__28133));
    InMux I__4629 (
            .O(N__28153),
            .I(N__28133));
    InMux I__4628 (
            .O(N__28152),
            .I(N__28108));
    InMux I__4627 (
            .O(N__28151),
            .I(N__28108));
    InMux I__4626 (
            .O(N__28150),
            .I(N__28108));
    InMux I__4625 (
            .O(N__28149),
            .I(N__28108));
    InMux I__4624 (
            .O(N__28148),
            .I(N__28108));
    InMux I__4623 (
            .O(N__28147),
            .I(N__28108));
    InMux I__4622 (
            .O(N__28146),
            .I(N__28103));
    InMux I__4621 (
            .O(N__28145),
            .I(N__28103));
    InMux I__4620 (
            .O(N__28144),
            .I(N__28098));
    LocalMux I__4619 (
            .O(N__28133),
            .I(N__28095));
    CascadeMux I__4618 (
            .O(N__28132),
            .I(N__28091));
    CascadeMux I__4617 (
            .O(N__28131),
            .I(N__28088));
    CascadeMux I__4616 (
            .O(N__28130),
            .I(N__28085));
    InMux I__4615 (
            .O(N__28129),
            .I(N__28074));
    InMux I__4614 (
            .O(N__28128),
            .I(N__28074));
    InMux I__4613 (
            .O(N__28127),
            .I(N__28074));
    InMux I__4612 (
            .O(N__28126),
            .I(N__28074));
    InMux I__4611 (
            .O(N__28125),
            .I(N__28063));
    InMux I__4610 (
            .O(N__28124),
            .I(N__28063));
    InMux I__4609 (
            .O(N__28123),
            .I(N__28063));
    InMux I__4608 (
            .O(N__28122),
            .I(N__28063));
    InMux I__4607 (
            .O(N__28121),
            .I(N__28063));
    LocalMux I__4606 (
            .O(N__28108),
            .I(N__28058));
    LocalMux I__4605 (
            .O(N__28103),
            .I(N__28058));
    InMux I__4604 (
            .O(N__28102),
            .I(N__28053));
    InMux I__4603 (
            .O(N__28101),
            .I(N__28053));
    LocalMux I__4602 (
            .O(N__28098),
            .I(N__28050));
    Span4Mux_v I__4601 (
            .O(N__28095),
            .I(N__28047));
    InMux I__4600 (
            .O(N__28094),
            .I(N__28044));
    InMux I__4599 (
            .O(N__28091),
            .I(N__28041));
    InMux I__4598 (
            .O(N__28088),
            .I(N__28032));
    InMux I__4597 (
            .O(N__28085),
            .I(N__28032));
    InMux I__4596 (
            .O(N__28084),
            .I(N__28032));
    InMux I__4595 (
            .O(N__28083),
            .I(N__28032));
    LocalMux I__4594 (
            .O(N__28074),
            .I(N__28025));
    LocalMux I__4593 (
            .O(N__28063),
            .I(N__28025));
    Span4Mux_v I__4592 (
            .O(N__28058),
            .I(N__28025));
    LocalMux I__4591 (
            .O(N__28053),
            .I(N__28018));
    Span4Mux_v I__4590 (
            .O(N__28050),
            .I(N__28018));
    Span4Mux_v I__4589 (
            .O(N__28047),
            .I(N__28018));
    LocalMux I__4588 (
            .O(N__28044),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    LocalMux I__4587 (
            .O(N__28041),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    LocalMux I__4586 (
            .O(N__28032),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__4585 (
            .O(N__28025),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__4584 (
            .O(N__28018),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    CascadeMux I__4583 (
            .O(N__28007),
            .I(N__27997));
    CascadeMux I__4582 (
            .O(N__28006),
            .I(N__27994));
    CascadeMux I__4581 (
            .O(N__28005),
            .I(N__27991));
    CascadeMux I__4580 (
            .O(N__28004),
            .I(N__27988));
    CascadeMux I__4579 (
            .O(N__28003),
            .I(N__27982));
    CascadeMux I__4578 (
            .O(N__28002),
            .I(N__27978));
    CascadeMux I__4577 (
            .O(N__28001),
            .I(N__27975));
    CascadeMux I__4576 (
            .O(N__28000),
            .I(N__27972));
    InMux I__4575 (
            .O(N__27997),
            .I(N__27959));
    InMux I__4574 (
            .O(N__27994),
            .I(N__27959));
    InMux I__4573 (
            .O(N__27991),
            .I(N__27948));
    InMux I__4572 (
            .O(N__27988),
            .I(N__27948));
    InMux I__4571 (
            .O(N__27987),
            .I(N__27948));
    InMux I__4570 (
            .O(N__27986),
            .I(N__27948));
    InMux I__4569 (
            .O(N__27985),
            .I(N__27948));
    InMux I__4568 (
            .O(N__27982),
            .I(N__27939));
    InMux I__4567 (
            .O(N__27981),
            .I(N__27939));
    InMux I__4566 (
            .O(N__27978),
            .I(N__27939));
    InMux I__4565 (
            .O(N__27975),
            .I(N__27939));
    InMux I__4564 (
            .O(N__27972),
            .I(N__27928));
    InMux I__4563 (
            .O(N__27971),
            .I(N__27928));
    InMux I__4562 (
            .O(N__27970),
            .I(N__27928));
    InMux I__4561 (
            .O(N__27969),
            .I(N__27928));
    InMux I__4560 (
            .O(N__27968),
            .I(N__27928));
    InMux I__4559 (
            .O(N__27967),
            .I(N__27923));
    InMux I__4558 (
            .O(N__27966),
            .I(N__27923));
    CascadeMux I__4557 (
            .O(N__27965),
            .I(N__27919));
    CascadeMux I__4556 (
            .O(N__27964),
            .I(N__27916));
    LocalMux I__4555 (
            .O(N__27959),
            .I(N__27907));
    LocalMux I__4554 (
            .O(N__27948),
            .I(N__27907));
    LocalMux I__4553 (
            .O(N__27939),
            .I(N__27907));
    LocalMux I__4552 (
            .O(N__27928),
            .I(N__27904));
    LocalMux I__4551 (
            .O(N__27923),
            .I(N__27900));
    InMux I__4550 (
            .O(N__27922),
            .I(N__27895));
    InMux I__4549 (
            .O(N__27919),
            .I(N__27895));
    InMux I__4548 (
            .O(N__27916),
            .I(N__27890));
    InMux I__4547 (
            .O(N__27915),
            .I(N__27890));
    CascadeMux I__4546 (
            .O(N__27914),
            .I(N__27887));
    Span4Mux_v I__4545 (
            .O(N__27907),
            .I(N__27874));
    Span4Mux_v I__4544 (
            .O(N__27904),
            .I(N__27874));
    InMux I__4543 (
            .O(N__27903),
            .I(N__27871));
    Span4Mux_v I__4542 (
            .O(N__27900),
            .I(N__27864));
    LocalMux I__4541 (
            .O(N__27895),
            .I(N__27864));
    LocalMux I__4540 (
            .O(N__27890),
            .I(N__27864));
    InMux I__4539 (
            .O(N__27887),
            .I(N__27861));
    InMux I__4538 (
            .O(N__27886),
            .I(N__27858));
    InMux I__4537 (
            .O(N__27885),
            .I(N__27855));
    CascadeMux I__4536 (
            .O(N__27884),
            .I(N__27852));
    CascadeMux I__4535 (
            .O(N__27883),
            .I(N__27849));
    CascadeMux I__4534 (
            .O(N__27882),
            .I(N__27846));
    CascadeMux I__4533 (
            .O(N__27881),
            .I(N__27843));
    CascadeMux I__4532 (
            .O(N__27880),
            .I(N__27840));
    InMux I__4531 (
            .O(N__27879),
            .I(N__27837));
    Span4Mux_h I__4530 (
            .O(N__27874),
            .I(N__27834));
    LocalMux I__4529 (
            .O(N__27871),
            .I(N__27831));
    Span4Mux_h I__4528 (
            .O(N__27864),
            .I(N__27828));
    LocalMux I__4527 (
            .O(N__27861),
            .I(N__27825));
    LocalMux I__4526 (
            .O(N__27858),
            .I(N__27820));
    LocalMux I__4525 (
            .O(N__27855),
            .I(N__27820));
    InMux I__4524 (
            .O(N__27852),
            .I(N__27813));
    InMux I__4523 (
            .O(N__27849),
            .I(N__27813));
    InMux I__4522 (
            .O(N__27846),
            .I(N__27813));
    InMux I__4521 (
            .O(N__27843),
            .I(N__27808));
    InMux I__4520 (
            .O(N__27840),
            .I(N__27808));
    LocalMux I__4519 (
            .O(N__27837),
            .I(N__27805));
    Sp12to4 I__4518 (
            .O(N__27834),
            .I(N__27802));
    Span4Mux_v I__4517 (
            .O(N__27831),
            .I(N__27793));
    Span4Mux_v I__4516 (
            .O(N__27828),
            .I(N__27793));
    Span4Mux_v I__4515 (
            .O(N__27825),
            .I(N__27793));
    Span4Mux_v I__4514 (
            .O(N__27820),
            .I(N__27793));
    LocalMux I__4513 (
            .O(N__27813),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__4512 (
            .O(N__27808),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4511 (
            .O(N__27805),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__4510 (
            .O(N__27802),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4509 (
            .O(N__27793),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__4508 (
            .O(N__27782),
            .I(N__27779));
    LocalMux I__4507 (
            .O(N__27779),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__4506 (
            .O(N__27776),
            .I(N__27773));
    InMux I__4505 (
            .O(N__27773),
            .I(N__27769));
    InMux I__4504 (
            .O(N__27772),
            .I(N__27766));
    LocalMux I__4503 (
            .O(N__27769),
            .I(N__27762));
    LocalMux I__4502 (
            .O(N__27766),
            .I(N__27759));
    InMux I__4501 (
            .O(N__27765),
            .I(N__27756));
    Span4Mux_h I__4500 (
            .O(N__27762),
            .I(N__27753));
    Span4Mux_v I__4499 (
            .O(N__27759),
            .I(N__27748));
    LocalMux I__4498 (
            .O(N__27756),
            .I(N__27748));
    Span4Mux_v I__4497 (
            .O(N__27753),
            .I(N__27744));
    Span4Mux_h I__4496 (
            .O(N__27748),
            .I(N__27741));
    InMux I__4495 (
            .O(N__27747),
            .I(N__27738));
    Odrv4 I__4494 (
            .O(N__27744),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__4493 (
            .O(N__27741),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__4492 (
            .O(N__27738),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__4491 (
            .O(N__27731),
            .I(N__27728));
    InMux I__4490 (
            .O(N__27728),
            .I(N__27725));
    LocalMux I__4489 (
            .O(N__27725),
            .I(N__27720));
    InMux I__4488 (
            .O(N__27724),
            .I(N__27717));
    InMux I__4487 (
            .O(N__27723),
            .I(N__27713));
    Span4Mux_h I__4486 (
            .O(N__27720),
            .I(N__27708));
    LocalMux I__4485 (
            .O(N__27717),
            .I(N__27708));
    InMux I__4484 (
            .O(N__27716),
            .I(N__27704));
    LocalMux I__4483 (
            .O(N__27713),
            .I(N__27701));
    Span4Mux_v I__4482 (
            .O(N__27708),
            .I(N__27698));
    InMux I__4481 (
            .O(N__27707),
            .I(N__27695));
    LocalMux I__4480 (
            .O(N__27704),
            .I(N__27692));
    Span4Mux_h I__4479 (
            .O(N__27701),
            .I(N__27689));
    Odrv4 I__4478 (
            .O(N__27698),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__4477 (
            .O(N__27695),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__4476 (
            .O(N__27692),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__4475 (
            .O(N__27689),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__4474 (
            .O(N__27680),
            .I(N__27677));
    LocalMux I__4473 (
            .O(N__27677),
            .I(N__27674));
    Odrv4 I__4472 (
            .O(N__27674),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    InMux I__4471 (
            .O(N__27671),
            .I(N__27668));
    LocalMux I__4470 (
            .O(N__27668),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ));
    InMux I__4469 (
            .O(N__27665),
            .I(N__27661));
    InMux I__4468 (
            .O(N__27664),
            .I(N__27658));
    LocalMux I__4467 (
            .O(N__27661),
            .I(N__27655));
    LocalMux I__4466 (
            .O(N__27658),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    Odrv4 I__4465 (
            .O(N__27655),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    InMux I__4464 (
            .O(N__27650),
            .I(N__27646));
    CascadeMux I__4463 (
            .O(N__27649),
            .I(N__27642));
    LocalMux I__4462 (
            .O(N__27646),
            .I(N__27638));
    CascadeMux I__4461 (
            .O(N__27645),
            .I(N__27635));
    InMux I__4460 (
            .O(N__27642),
            .I(N__27630));
    InMux I__4459 (
            .O(N__27641),
            .I(N__27630));
    Span4Mux_h I__4458 (
            .O(N__27638),
            .I(N__27626));
    InMux I__4457 (
            .O(N__27635),
            .I(N__27623));
    LocalMux I__4456 (
            .O(N__27630),
            .I(N__27620));
    InMux I__4455 (
            .O(N__27629),
            .I(N__27617));
    Odrv4 I__4454 (
            .O(N__27626),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__4453 (
            .O(N__27623),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__4452 (
            .O(N__27620),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__4451 (
            .O(N__27617),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    CascadeMux I__4450 (
            .O(N__27608),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_ ));
    InMux I__4449 (
            .O(N__27605),
            .I(N__27602));
    LocalMux I__4448 (
            .O(N__27602),
            .I(N__27599));
    Odrv4 I__4447 (
            .O(N__27599),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    InMux I__4446 (
            .O(N__27596),
            .I(N__27593));
    LocalMux I__4445 (
            .O(N__27593),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ));
    InMux I__4444 (
            .O(N__27590),
            .I(N__27586));
    InMux I__4443 (
            .O(N__27589),
            .I(N__27583));
    LocalMux I__4442 (
            .O(N__27586),
            .I(N__27580));
    LocalMux I__4441 (
            .O(N__27583),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    Odrv12 I__4440 (
            .O(N__27580),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    CascadeMux I__4439 (
            .O(N__27575),
            .I(N__27571));
    CascadeMux I__4438 (
            .O(N__27574),
            .I(N__27568));
    InMux I__4437 (
            .O(N__27571),
            .I(N__27564));
    InMux I__4436 (
            .O(N__27568),
            .I(N__27561));
    InMux I__4435 (
            .O(N__27567),
            .I(N__27557));
    LocalMux I__4434 (
            .O(N__27564),
            .I(N__27554));
    LocalMux I__4433 (
            .O(N__27561),
            .I(N__27551));
    InMux I__4432 (
            .O(N__27560),
            .I(N__27547));
    LocalMux I__4431 (
            .O(N__27557),
            .I(N__27544));
    Span4Mux_h I__4430 (
            .O(N__27554),
            .I(N__27541));
    Span4Mux_v I__4429 (
            .O(N__27551),
            .I(N__27538));
    InMux I__4428 (
            .O(N__27550),
            .I(N__27535));
    LocalMux I__4427 (
            .O(N__27547),
            .I(N__27532));
    Span4Mux_v I__4426 (
            .O(N__27544),
            .I(N__27529));
    Odrv4 I__4425 (
            .O(N__27541),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__4424 (
            .O(N__27538),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__4423 (
            .O(N__27535),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__4422 (
            .O(N__27532),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__4421 (
            .O(N__27529),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__4420 (
            .O(N__27518),
            .I(N__27515));
    LocalMux I__4419 (
            .O(N__27515),
            .I(N__27512));
    Odrv4 I__4418 (
            .O(N__27512),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__4417 (
            .O(N__27509),
            .I(N__27506));
    LocalMux I__4416 (
            .O(N__27506),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ));
    InMux I__4415 (
            .O(N__27503),
            .I(N__27500));
    LocalMux I__4414 (
            .O(N__27500),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__4413 (
            .O(N__27497),
            .I(N__27494));
    LocalMux I__4412 (
            .O(N__27494),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ));
    InMux I__4411 (
            .O(N__27491),
            .I(N__27488));
    LocalMux I__4410 (
            .O(N__27488),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__4409 (
            .O(N__27485),
            .I(N__27482));
    LocalMux I__4408 (
            .O(N__27482),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ));
    CascadeMux I__4407 (
            .O(N__27479),
            .I(N__27476));
    InMux I__4406 (
            .O(N__27476),
            .I(N__27473));
    LocalMux I__4405 (
            .O(N__27473),
            .I(N__27470));
    Odrv4 I__4404 (
            .O(N__27470),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__4403 (
            .O(N__27467),
            .I(N__27464));
    LocalMux I__4402 (
            .O(N__27464),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ));
    CascadeMux I__4401 (
            .O(N__27461),
            .I(N__27458));
    InMux I__4400 (
            .O(N__27458),
            .I(N__27454));
    InMux I__4399 (
            .O(N__27457),
            .I(N__27450));
    LocalMux I__4398 (
            .O(N__27454),
            .I(N__27447));
    InMux I__4397 (
            .O(N__27453),
            .I(N__27444));
    LocalMux I__4396 (
            .O(N__27450),
            .I(N__27439));
    Span4Mux_h I__4395 (
            .O(N__27447),
            .I(N__27436));
    LocalMux I__4394 (
            .O(N__27444),
            .I(N__27433));
    InMux I__4393 (
            .O(N__27443),
            .I(N__27428));
    InMux I__4392 (
            .O(N__27442),
            .I(N__27428));
    Odrv4 I__4391 (
            .O(N__27439),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__4390 (
            .O(N__27436),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__4389 (
            .O(N__27433),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__4388 (
            .O(N__27428),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__4387 (
            .O(N__27419),
            .I(N__27416));
    LocalMux I__4386 (
            .O(N__27416),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    InMux I__4385 (
            .O(N__27413),
            .I(N__27410));
    LocalMux I__4384 (
            .O(N__27410),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ));
    CascadeMux I__4383 (
            .O(N__27407),
            .I(N__27403));
    InMux I__4382 (
            .O(N__27406),
            .I(N__27398));
    InMux I__4381 (
            .O(N__27403),
            .I(N__27395));
    InMux I__4380 (
            .O(N__27402),
            .I(N__27392));
    InMux I__4379 (
            .O(N__27401),
            .I(N__27388));
    LocalMux I__4378 (
            .O(N__27398),
            .I(N__27385));
    LocalMux I__4377 (
            .O(N__27395),
            .I(N__27382));
    LocalMux I__4376 (
            .O(N__27392),
            .I(N__27379));
    InMux I__4375 (
            .O(N__27391),
            .I(N__27376));
    LocalMux I__4374 (
            .O(N__27388),
            .I(N__27373));
    Span4Mux_h I__4373 (
            .O(N__27385),
            .I(N__27370));
    Odrv4 I__4372 (
            .O(N__27382),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4371 (
            .O(N__27379),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__4370 (
            .O(N__27376),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv12 I__4369 (
            .O(N__27373),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4368 (
            .O(N__27370),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__4367 (
            .O(N__27359),
            .I(N__27356));
    LocalMux I__4366 (
            .O(N__27356),
            .I(N__27353));
    Odrv4 I__4365 (
            .O(N__27353),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    InMux I__4364 (
            .O(N__27350),
            .I(N__27347));
    LocalMux I__4363 (
            .O(N__27347),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ));
    InMux I__4362 (
            .O(N__27344),
            .I(N__27341));
    LocalMux I__4361 (
            .O(N__27341),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    InMux I__4360 (
            .O(N__27338),
            .I(N__27335));
    LocalMux I__4359 (
            .O(N__27335),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ));
    InMux I__4358 (
            .O(N__27332),
            .I(N__27329));
    LocalMux I__4357 (
            .O(N__27329),
            .I(N__27326));
    Odrv12 I__4356 (
            .O(N__27326),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    CascadeMux I__4355 (
            .O(N__27323),
            .I(N__27320));
    InMux I__4354 (
            .O(N__27320),
            .I(N__27317));
    LocalMux I__4353 (
            .O(N__27317),
            .I(N__27314));
    Odrv4 I__4352 (
            .O(N__27314),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ));
    InMux I__4351 (
            .O(N__27311),
            .I(N__27308));
    LocalMux I__4350 (
            .O(N__27308),
            .I(N__27305));
    Odrv4 I__4349 (
            .O(N__27305),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__4348 (
            .O(N__27302),
            .I(N__27298));
    InMux I__4347 (
            .O(N__27301),
            .I(N__27294));
    LocalMux I__4346 (
            .O(N__27298),
            .I(N__27290));
    InMux I__4345 (
            .O(N__27297),
            .I(N__27287));
    LocalMux I__4344 (
            .O(N__27294),
            .I(N__27284));
    CascadeMux I__4343 (
            .O(N__27293),
            .I(N__27281));
    Span4Mux_v I__4342 (
            .O(N__27290),
            .I(N__27276));
    LocalMux I__4341 (
            .O(N__27287),
            .I(N__27276));
    Span4Mux_h I__4340 (
            .O(N__27284),
            .I(N__27272));
    InMux I__4339 (
            .O(N__27281),
            .I(N__27269));
    Span4Mux_h I__4338 (
            .O(N__27276),
            .I(N__27266));
    InMux I__4337 (
            .O(N__27275),
            .I(N__27263));
    Span4Mux_v I__4336 (
            .O(N__27272),
            .I(N__27260));
    LocalMux I__4335 (
            .O(N__27269),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4334 (
            .O(N__27266),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4333 (
            .O(N__27263),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4332 (
            .O(N__27260),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__4331 (
            .O(N__27251),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__4330 (
            .O(N__27248),
            .I(bfn_11_11_0_));
    InMux I__4329 (
            .O(N__27245),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__4328 (
            .O(N__27242),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__4327 (
            .O(N__27239),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__4326 (
            .O(N__27236),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__4325 (
            .O(N__27233),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__4324 (
            .O(N__27230),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__4323 (
            .O(N__27227),
            .I(N__27223));
    CascadeMux I__4322 (
            .O(N__27226),
            .I(N__27220));
    LocalMux I__4321 (
            .O(N__27223),
            .I(N__27215));
    InMux I__4320 (
            .O(N__27220),
            .I(N__27212));
    InMux I__4319 (
            .O(N__27219),
            .I(N__27209));
    CascadeMux I__4318 (
            .O(N__27218),
            .I(N__27205));
    Span4Mux_v I__4317 (
            .O(N__27215),
            .I(N__27200));
    LocalMux I__4316 (
            .O(N__27212),
            .I(N__27200));
    LocalMux I__4315 (
            .O(N__27209),
            .I(N__27197));
    InMux I__4314 (
            .O(N__27208),
            .I(N__27192));
    InMux I__4313 (
            .O(N__27205),
            .I(N__27192));
    Odrv4 I__4312 (
            .O(N__27200),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__4311 (
            .O(N__27197),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__4310 (
            .O(N__27192),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__4309 (
            .O(N__27185),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    InMux I__4308 (
            .O(N__27182),
            .I(N__27179));
    LocalMux I__4307 (
            .O(N__27179),
            .I(N__27176));
    Odrv4 I__4306 (
            .O(N__27176),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ));
    InMux I__4305 (
            .O(N__27173),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    InMux I__4304 (
            .O(N__27170),
            .I(N__27167));
    LocalMux I__4303 (
            .O(N__27167),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    InMux I__4302 (
            .O(N__27164),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__4301 (
            .O(N__27161),
            .I(bfn_11_10_0_));
    InMux I__4300 (
            .O(N__27158),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__4299 (
            .O(N__27155),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__4298 (
            .O(N__27152),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__4297 (
            .O(N__27149),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__4296 (
            .O(N__27146),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__4295 (
            .O(N__27143),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__4294 (
            .O(N__27140),
            .I(N__27137));
    LocalMux I__4293 (
            .O(N__27137),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    InMux I__4292 (
            .O(N__27134),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__4291 (
            .O(N__27131),
            .I(N__27128));
    LocalMux I__4290 (
            .O(N__27128),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__4289 (
            .O(N__27125),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    InMux I__4288 (
            .O(N__27122),
            .I(N__27119));
    LocalMux I__4287 (
            .O(N__27119),
            .I(N__27116));
    Odrv12 I__4286 (
            .O(N__27116),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__4285 (
            .O(N__27113),
            .I(N__27110));
    LocalMux I__4284 (
            .O(N__27110),
            .I(N__27107));
    Odrv4 I__4283 (
            .O(N__27107),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__4282 (
            .O(N__27104),
            .I(bfn_11_9_0_));
    InMux I__4281 (
            .O(N__27101),
            .I(N__27098));
    LocalMux I__4280 (
            .O(N__27098),
            .I(N__27095));
    Odrv12 I__4279 (
            .O(N__27095),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__4278 (
            .O(N__27092),
            .I(N__27089));
    LocalMux I__4277 (
            .O(N__27089),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__4276 (
            .O(N__27086),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    InMux I__4275 (
            .O(N__27083),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__4274 (
            .O(N__27080),
            .I(N__27077));
    LocalMux I__4273 (
            .O(N__27077),
            .I(N__27074));
    Span4Mux_v I__4272 (
            .O(N__27074),
            .I(N__27071));
    Odrv4 I__4271 (
            .O(N__27071),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__4270 (
            .O(N__27068),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__4269 (
            .O(N__27065),
            .I(N__27062));
    LocalMux I__4268 (
            .O(N__27062),
            .I(N__27059));
    Odrv4 I__4267 (
            .O(N__27059),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ));
    InMux I__4266 (
            .O(N__27056),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__4265 (
            .O(N__27053),
            .I(N__27050));
    LocalMux I__4264 (
            .O(N__27050),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ));
    InMux I__4263 (
            .O(N__27047),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__4262 (
            .O(N__27044),
            .I(N__27041));
    LocalMux I__4261 (
            .O(N__27041),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    InMux I__4260 (
            .O(N__27038),
            .I(N__27035));
    LocalMux I__4259 (
            .O(N__27035),
            .I(N__27032));
    Odrv4 I__4258 (
            .O(N__27032),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    CascadeMux I__4257 (
            .O(N__27029),
            .I(N__27026));
    InMux I__4256 (
            .O(N__27026),
            .I(N__27023));
    LocalMux I__4255 (
            .O(N__27023),
            .I(N__27020));
    Odrv4 I__4254 (
            .O(N__27020),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__4253 (
            .O(N__27017),
            .I(N__27014));
    LocalMux I__4252 (
            .O(N__27014),
            .I(N__27011));
    Span4Mux_v I__4251 (
            .O(N__27011),
            .I(N__27007));
    InMux I__4250 (
            .O(N__27010),
            .I(N__27004));
    Odrv4 I__4249 (
            .O(N__27007),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    LocalMux I__4248 (
            .O(N__27004),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__4247 (
            .O(N__26999),
            .I(N__26996));
    LocalMux I__4246 (
            .O(N__26996),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__4245 (
            .O(N__26993),
            .I(N__26990));
    LocalMux I__4244 (
            .O(N__26990),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__4243 (
            .O(N__26987),
            .I(N__26984));
    LocalMux I__4242 (
            .O(N__26984),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__4241 (
            .O(N__26981),
            .I(N__26978));
    LocalMux I__4240 (
            .O(N__26978),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__4239 (
            .O(N__26975),
            .I(N__26972));
    LocalMux I__4238 (
            .O(N__26972),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__4237 (
            .O(N__26969),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    InMux I__4236 (
            .O(N__26966),
            .I(N__26963));
    LocalMux I__4235 (
            .O(N__26963),
            .I(N__26960));
    Odrv4 I__4234 (
            .O(N__26960),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__4233 (
            .O(N__26957),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    CascadeMux I__4232 (
            .O(N__26954),
            .I(N__26951));
    InMux I__4231 (
            .O(N__26951),
            .I(N__26948));
    LocalMux I__4230 (
            .O(N__26948),
            .I(N__26945));
    Span4Mux_v I__4229 (
            .O(N__26945),
            .I(N__26942));
    Odrv4 I__4228 (
            .O(N__26942),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    InMux I__4227 (
            .O(N__26939),
            .I(N__26901));
    InMux I__4226 (
            .O(N__26938),
            .I(N__26901));
    InMux I__4225 (
            .O(N__26937),
            .I(N__26901));
    InMux I__4224 (
            .O(N__26936),
            .I(N__26901));
    InMux I__4223 (
            .O(N__26935),
            .I(N__26892));
    InMux I__4222 (
            .O(N__26934),
            .I(N__26892));
    InMux I__4221 (
            .O(N__26933),
            .I(N__26892));
    InMux I__4220 (
            .O(N__26932),
            .I(N__26892));
    InMux I__4219 (
            .O(N__26931),
            .I(N__26883));
    InMux I__4218 (
            .O(N__26930),
            .I(N__26883));
    InMux I__4217 (
            .O(N__26929),
            .I(N__26883));
    InMux I__4216 (
            .O(N__26928),
            .I(N__26883));
    InMux I__4215 (
            .O(N__26927),
            .I(N__26874));
    InMux I__4214 (
            .O(N__26926),
            .I(N__26874));
    InMux I__4213 (
            .O(N__26925),
            .I(N__26874));
    InMux I__4212 (
            .O(N__26924),
            .I(N__26874));
    InMux I__4211 (
            .O(N__26923),
            .I(N__26869));
    InMux I__4210 (
            .O(N__26922),
            .I(N__26869));
    InMux I__4209 (
            .O(N__26921),
            .I(N__26860));
    InMux I__4208 (
            .O(N__26920),
            .I(N__26860));
    InMux I__4207 (
            .O(N__26919),
            .I(N__26860));
    InMux I__4206 (
            .O(N__26918),
            .I(N__26860));
    InMux I__4205 (
            .O(N__26917),
            .I(N__26851));
    InMux I__4204 (
            .O(N__26916),
            .I(N__26851));
    InMux I__4203 (
            .O(N__26915),
            .I(N__26851));
    InMux I__4202 (
            .O(N__26914),
            .I(N__26851));
    InMux I__4201 (
            .O(N__26913),
            .I(N__26842));
    InMux I__4200 (
            .O(N__26912),
            .I(N__26842));
    InMux I__4199 (
            .O(N__26911),
            .I(N__26842));
    InMux I__4198 (
            .O(N__26910),
            .I(N__26842));
    LocalMux I__4197 (
            .O(N__26901),
            .I(N__26839));
    LocalMux I__4196 (
            .O(N__26892),
            .I(N__26836));
    LocalMux I__4195 (
            .O(N__26883),
            .I(N__26831));
    LocalMux I__4194 (
            .O(N__26874),
            .I(N__26831));
    LocalMux I__4193 (
            .O(N__26869),
            .I(N__26828));
    LocalMux I__4192 (
            .O(N__26860),
            .I(N__26825));
    LocalMux I__4191 (
            .O(N__26851),
            .I(N__26820));
    LocalMux I__4190 (
            .O(N__26842),
            .I(N__26820));
    Span4Mux_h I__4189 (
            .O(N__26839),
            .I(N__26817));
    Span4Mux_h I__4188 (
            .O(N__26836),
            .I(N__26814));
    Span4Mux_h I__4187 (
            .O(N__26831),
            .I(N__26811));
    Span4Mux_v I__4186 (
            .O(N__26828),
            .I(N__26806));
    Span4Mux_v I__4185 (
            .O(N__26825),
            .I(N__26806));
    Span4Mux_h I__4184 (
            .O(N__26820),
            .I(N__26803));
    Span4Mux_v I__4183 (
            .O(N__26817),
            .I(N__26798));
    Span4Mux_v I__4182 (
            .O(N__26814),
            .I(N__26798));
    Span4Mux_v I__4181 (
            .O(N__26811),
            .I(N__26795));
    Odrv4 I__4180 (
            .O(N__26806),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__4179 (
            .O(N__26803),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__4178 (
            .O(N__26798),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__4177 (
            .O(N__26795),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__4176 (
            .O(N__26786),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CascadeMux I__4175 (
            .O(N__26783),
            .I(N__26780));
    InMux I__4174 (
            .O(N__26780),
            .I(N__26776));
    InMux I__4173 (
            .O(N__26779),
            .I(N__26773));
    LocalMux I__4172 (
            .O(N__26776),
            .I(N__26770));
    LocalMux I__4171 (
            .O(N__26773),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__4170 (
            .O(N__26770),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    InMux I__4169 (
            .O(N__26765),
            .I(N__26759));
    InMux I__4168 (
            .O(N__26764),
            .I(N__26756));
    InMux I__4167 (
            .O(N__26763),
            .I(N__26751));
    InMux I__4166 (
            .O(N__26762),
            .I(N__26751));
    LocalMux I__4165 (
            .O(N__26759),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__4164 (
            .O(N__26756),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__4163 (
            .O(N__26751),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    CascadeMux I__4162 (
            .O(N__26744),
            .I(\delay_measurement_inst.N_39_cascade_ ));
    InMux I__4161 (
            .O(N__26741),
            .I(N__26738));
    LocalMux I__4160 (
            .O(N__26738),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__4159 (
            .O(N__26735),
            .I(N__26732));
    LocalMux I__4158 (
            .O(N__26732),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    CascadeMux I__4157 (
            .O(N__26729),
            .I(N__26726));
    InMux I__4156 (
            .O(N__26726),
            .I(N__26723));
    LocalMux I__4155 (
            .O(N__26723),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_26 ));
    InMux I__4154 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__4153 (
            .O(N__26717),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__4152 (
            .O(N__26714),
            .I(N__26711));
    LocalMux I__4151 (
            .O(N__26711),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__4150 (
            .O(N__26708),
            .I(N__26705));
    LocalMux I__4149 (
            .O(N__26705),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__4148 (
            .O(N__26702),
            .I(N__26699));
    LocalMux I__4147 (
            .O(N__26699),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ));
    CascadeMux I__4146 (
            .O(N__26696),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ));
    InMux I__4145 (
            .O(N__26693),
            .I(N__26690));
    LocalMux I__4144 (
            .O(N__26690),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ));
    InMux I__4143 (
            .O(N__26687),
            .I(N__26684));
    LocalMux I__4142 (
            .O(N__26684),
            .I(N__26681));
    Span4Mux_h I__4141 (
            .O(N__26681),
            .I(N__26677));
    InMux I__4140 (
            .O(N__26680),
            .I(N__26674));
    Odrv4 I__4139 (
            .O(N__26677),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    LocalMux I__4138 (
            .O(N__26674),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    InMux I__4137 (
            .O(N__26669),
            .I(N__26665));
    InMux I__4136 (
            .O(N__26668),
            .I(N__26662));
    LocalMux I__4135 (
            .O(N__26665),
            .I(\delay_measurement_inst.elapsed_time_hc_27 ));
    LocalMux I__4134 (
            .O(N__26662),
            .I(\delay_measurement_inst.elapsed_time_hc_27 ));
    IoInMux I__4133 (
            .O(N__26657),
            .I(N__26654));
    LocalMux I__4132 (
            .O(N__26654),
            .I(N__26651));
    Span4Mux_s3_v I__4131 (
            .O(N__26651),
            .I(N__26648));
    Sp12to4 I__4130 (
            .O(N__26648),
            .I(N__26645));
    Odrv12 I__4129 (
            .O(N__26645),
            .I(s3_phy_c));
    CascadeMux I__4128 (
            .O(N__26642),
            .I(N__26638));
    CascadeMux I__4127 (
            .O(N__26641),
            .I(N__26635));
    InMux I__4126 (
            .O(N__26638),
            .I(N__26629));
    InMux I__4125 (
            .O(N__26635),
            .I(N__26629));
    InMux I__4124 (
            .O(N__26634),
            .I(N__26626));
    LocalMux I__4123 (
            .O(N__26629),
            .I(N__26623));
    LocalMux I__4122 (
            .O(N__26626),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__4121 (
            .O(N__26623),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__4120 (
            .O(N__26618),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__4119 (
            .O(N__26615),
            .I(N__26612));
    InMux I__4118 (
            .O(N__26612),
            .I(N__26608));
    InMux I__4117 (
            .O(N__26611),
            .I(N__26604));
    LocalMux I__4116 (
            .O(N__26608),
            .I(N__26601));
    InMux I__4115 (
            .O(N__26607),
            .I(N__26598));
    LocalMux I__4114 (
            .O(N__26604),
            .I(N__26593));
    Span4Mux_h I__4113 (
            .O(N__26601),
            .I(N__26593));
    LocalMux I__4112 (
            .O(N__26598),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__4111 (
            .O(N__26593),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__4110 (
            .O(N__26588),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__4109 (
            .O(N__26585),
            .I(N__26579));
    InMux I__4108 (
            .O(N__26584),
            .I(N__26579));
    LocalMux I__4107 (
            .O(N__26579),
            .I(N__26575));
    InMux I__4106 (
            .O(N__26578),
            .I(N__26572));
    Span4Mux_h I__4105 (
            .O(N__26575),
            .I(N__26569));
    LocalMux I__4104 (
            .O(N__26572),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__4103 (
            .O(N__26569),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__4102 (
            .O(N__26564),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__4101 (
            .O(N__26561),
            .I(N__26558));
    InMux I__4100 (
            .O(N__26558),
            .I(N__26554));
    CascadeMux I__4099 (
            .O(N__26557),
            .I(N__26550));
    LocalMux I__4098 (
            .O(N__26554),
            .I(N__26547));
    InMux I__4097 (
            .O(N__26553),
            .I(N__26544));
    InMux I__4096 (
            .O(N__26550),
            .I(N__26541));
    Odrv4 I__4095 (
            .O(N__26547),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__4094 (
            .O(N__26544),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__4093 (
            .O(N__26541),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__4092 (
            .O(N__26534),
            .I(bfn_10_20_0_));
    CascadeMux I__4091 (
            .O(N__26531),
            .I(N__26528));
    InMux I__4090 (
            .O(N__26528),
            .I(N__26525));
    LocalMux I__4089 (
            .O(N__26525),
            .I(N__26520));
    CascadeMux I__4088 (
            .O(N__26524),
            .I(N__26517));
    InMux I__4087 (
            .O(N__26523),
            .I(N__26514));
    Span4Mux_h I__4086 (
            .O(N__26520),
            .I(N__26511));
    InMux I__4085 (
            .O(N__26517),
            .I(N__26508));
    LocalMux I__4084 (
            .O(N__26514),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__4083 (
            .O(N__26511),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__4082 (
            .O(N__26508),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__4081 (
            .O(N__26501),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__4080 (
            .O(N__26498),
            .I(N__26495));
    InMux I__4079 (
            .O(N__26495),
            .I(N__26491));
    InMux I__4078 (
            .O(N__26494),
            .I(N__26488));
    LocalMux I__4077 (
            .O(N__26491),
            .I(N__26482));
    LocalMux I__4076 (
            .O(N__26488),
            .I(N__26482));
    InMux I__4075 (
            .O(N__26487),
            .I(N__26479));
    Span4Mux_v I__4074 (
            .O(N__26482),
            .I(N__26476));
    LocalMux I__4073 (
            .O(N__26479),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__4072 (
            .O(N__26476),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__4071 (
            .O(N__26471),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__4070 (
            .O(N__26468),
            .I(N__26461));
    InMux I__4069 (
            .O(N__26467),
            .I(N__26461));
    InMux I__4068 (
            .O(N__26466),
            .I(N__26458));
    LocalMux I__4067 (
            .O(N__26461),
            .I(N__26455));
    LocalMux I__4066 (
            .O(N__26458),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__4065 (
            .O(N__26455),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__4064 (
            .O(N__26450),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__4063 (
            .O(N__26447),
            .I(N__26443));
    InMux I__4062 (
            .O(N__26446),
            .I(N__26440));
    LocalMux I__4061 (
            .O(N__26443),
            .I(N__26437));
    LocalMux I__4060 (
            .O(N__26440),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__4059 (
            .O(N__26437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__4058 (
            .O(N__26432),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__4057 (
            .O(N__26429),
            .I(N__26422));
    InMux I__4056 (
            .O(N__26428),
            .I(N__26422));
    InMux I__4055 (
            .O(N__26427),
            .I(N__26419));
    LocalMux I__4054 (
            .O(N__26422),
            .I(N__26416));
    LocalMux I__4053 (
            .O(N__26419),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__4052 (
            .O(N__26416),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__4051 (
            .O(N__26411),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__4050 (
            .O(N__26408),
            .I(N__26404));
    CascadeMux I__4049 (
            .O(N__26407),
            .I(N__26401));
    InMux I__4048 (
            .O(N__26404),
            .I(N__26395));
    InMux I__4047 (
            .O(N__26401),
            .I(N__26395));
    InMux I__4046 (
            .O(N__26400),
            .I(N__26392));
    LocalMux I__4045 (
            .O(N__26395),
            .I(N__26389));
    LocalMux I__4044 (
            .O(N__26392),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__4043 (
            .O(N__26389),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__4042 (
            .O(N__26384),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__4041 (
            .O(N__26381),
            .I(N__26378));
    InMux I__4040 (
            .O(N__26378),
            .I(N__26374));
    InMux I__4039 (
            .O(N__26377),
            .I(N__26370));
    LocalMux I__4038 (
            .O(N__26374),
            .I(N__26367));
    InMux I__4037 (
            .O(N__26373),
            .I(N__26364));
    LocalMux I__4036 (
            .O(N__26370),
            .I(N__26359));
    Span4Mux_h I__4035 (
            .O(N__26367),
            .I(N__26359));
    LocalMux I__4034 (
            .O(N__26364),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__4033 (
            .O(N__26359),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__4032 (
            .O(N__26354),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__4031 (
            .O(N__26351),
            .I(N__26345));
    InMux I__4030 (
            .O(N__26350),
            .I(N__26345));
    LocalMux I__4029 (
            .O(N__26345),
            .I(N__26341));
    InMux I__4028 (
            .O(N__26344),
            .I(N__26338));
    Span4Mux_h I__4027 (
            .O(N__26341),
            .I(N__26335));
    LocalMux I__4026 (
            .O(N__26338),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__4025 (
            .O(N__26335),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__4024 (
            .O(N__26330),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__4023 (
            .O(N__26327),
            .I(N__26323));
    CascadeMux I__4022 (
            .O(N__26326),
            .I(N__26319));
    LocalMux I__4021 (
            .O(N__26323),
            .I(N__26316));
    InMux I__4020 (
            .O(N__26322),
            .I(N__26313));
    InMux I__4019 (
            .O(N__26319),
            .I(N__26310));
    Span4Mux_h I__4018 (
            .O(N__26316),
            .I(N__26307));
    LocalMux I__4017 (
            .O(N__26313),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__4016 (
            .O(N__26310),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__4015 (
            .O(N__26307),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__4014 (
            .O(N__26300),
            .I(bfn_10_19_0_));
    CascadeMux I__4013 (
            .O(N__26297),
            .I(N__26294));
    InMux I__4012 (
            .O(N__26294),
            .I(N__26291));
    LocalMux I__4011 (
            .O(N__26291),
            .I(N__26286));
    CascadeMux I__4010 (
            .O(N__26290),
            .I(N__26283));
    InMux I__4009 (
            .O(N__26289),
            .I(N__26280));
    Span4Mux_h I__4008 (
            .O(N__26286),
            .I(N__26277));
    InMux I__4007 (
            .O(N__26283),
            .I(N__26274));
    LocalMux I__4006 (
            .O(N__26280),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__4005 (
            .O(N__26277),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__4004 (
            .O(N__26274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__4003 (
            .O(N__26267),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__4002 (
            .O(N__26264),
            .I(N__26260));
    CascadeMux I__4001 (
            .O(N__26263),
            .I(N__26257));
    InMux I__4000 (
            .O(N__26260),
            .I(N__26251));
    InMux I__3999 (
            .O(N__26257),
            .I(N__26251));
    InMux I__3998 (
            .O(N__26256),
            .I(N__26248));
    LocalMux I__3997 (
            .O(N__26251),
            .I(N__26245));
    LocalMux I__3996 (
            .O(N__26248),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__3995 (
            .O(N__26245),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__3994 (
            .O(N__26240),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__3993 (
            .O(N__26237),
            .I(N__26230));
    InMux I__3992 (
            .O(N__26236),
            .I(N__26230));
    InMux I__3991 (
            .O(N__26235),
            .I(N__26227));
    LocalMux I__3990 (
            .O(N__26230),
            .I(N__26224));
    LocalMux I__3989 (
            .O(N__26227),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__3988 (
            .O(N__26224),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__3987 (
            .O(N__26219),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__3986 (
            .O(N__26216),
            .I(N__26209));
    InMux I__3985 (
            .O(N__26215),
            .I(N__26209));
    InMux I__3984 (
            .O(N__26214),
            .I(N__26206));
    LocalMux I__3983 (
            .O(N__26209),
            .I(N__26203));
    LocalMux I__3982 (
            .O(N__26206),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__3981 (
            .O(N__26203),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__3980 (
            .O(N__26198),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__3979 (
            .O(N__26195),
            .I(N__26191));
    CascadeMux I__3978 (
            .O(N__26194),
            .I(N__26188));
    InMux I__3977 (
            .O(N__26191),
            .I(N__26183));
    InMux I__3976 (
            .O(N__26188),
            .I(N__26183));
    LocalMux I__3975 (
            .O(N__26183),
            .I(N__26179));
    InMux I__3974 (
            .O(N__26182),
            .I(N__26176));
    Span4Mux_h I__3973 (
            .O(N__26179),
            .I(N__26173));
    LocalMux I__3972 (
            .O(N__26176),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__3971 (
            .O(N__26173),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__3970 (
            .O(N__26168),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__3969 (
            .O(N__26165),
            .I(N__26161));
    CascadeMux I__3968 (
            .O(N__26164),
            .I(N__26158));
    InMux I__3967 (
            .O(N__26161),
            .I(N__26152));
    InMux I__3966 (
            .O(N__26158),
            .I(N__26152));
    InMux I__3965 (
            .O(N__26157),
            .I(N__26149));
    LocalMux I__3964 (
            .O(N__26152),
            .I(N__26146));
    LocalMux I__3963 (
            .O(N__26149),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__3962 (
            .O(N__26146),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__3961 (
            .O(N__26141),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__3960 (
            .O(N__26138),
            .I(N__26131));
    InMux I__3959 (
            .O(N__26137),
            .I(N__26131));
    InMux I__3958 (
            .O(N__26136),
            .I(N__26128));
    LocalMux I__3957 (
            .O(N__26131),
            .I(N__26125));
    LocalMux I__3956 (
            .O(N__26128),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__3955 (
            .O(N__26125),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__3954 (
            .O(N__26120),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__3953 (
            .O(N__26117),
            .I(N__26111));
    InMux I__3952 (
            .O(N__26116),
            .I(N__26111));
    LocalMux I__3951 (
            .O(N__26111),
            .I(N__26107));
    InMux I__3950 (
            .O(N__26110),
            .I(N__26104));
    Span4Mux_h I__3949 (
            .O(N__26107),
            .I(N__26101));
    LocalMux I__3948 (
            .O(N__26104),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__3947 (
            .O(N__26101),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__3946 (
            .O(N__26096),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__3945 (
            .O(N__26093),
            .I(N__26090));
    LocalMux I__3944 (
            .O(N__26090),
            .I(N__26086));
    CascadeMux I__3943 (
            .O(N__26089),
            .I(N__26082));
    Span4Mux_v I__3942 (
            .O(N__26086),
            .I(N__26079));
    InMux I__3941 (
            .O(N__26085),
            .I(N__26076));
    InMux I__3940 (
            .O(N__26082),
            .I(N__26073));
    Odrv4 I__3939 (
            .O(N__26079),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__3938 (
            .O(N__26076),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__3937 (
            .O(N__26073),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__3936 (
            .O(N__26066),
            .I(bfn_10_18_0_));
    CascadeMux I__3935 (
            .O(N__26063),
            .I(N__26060));
    InMux I__3934 (
            .O(N__26060),
            .I(N__26057));
    LocalMux I__3933 (
            .O(N__26057),
            .I(N__26052));
    CascadeMux I__3932 (
            .O(N__26056),
            .I(N__26049));
    InMux I__3931 (
            .O(N__26055),
            .I(N__26046));
    Span4Mux_h I__3930 (
            .O(N__26052),
            .I(N__26043));
    InMux I__3929 (
            .O(N__26049),
            .I(N__26040));
    LocalMux I__3928 (
            .O(N__26046),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__3927 (
            .O(N__26043),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__3926 (
            .O(N__26040),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__3925 (
            .O(N__26033),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__3924 (
            .O(N__26030),
            .I(N__26026));
    CascadeMux I__3923 (
            .O(N__26029),
            .I(N__26023));
    InMux I__3922 (
            .O(N__26026),
            .I(N__26017));
    InMux I__3921 (
            .O(N__26023),
            .I(N__26017));
    InMux I__3920 (
            .O(N__26022),
            .I(N__26014));
    LocalMux I__3919 (
            .O(N__26017),
            .I(N__26011));
    LocalMux I__3918 (
            .O(N__26014),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__3917 (
            .O(N__26011),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__3916 (
            .O(N__26006),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__3915 (
            .O(N__26003),
            .I(N__25996));
    InMux I__3914 (
            .O(N__26002),
            .I(N__25996));
    InMux I__3913 (
            .O(N__26001),
            .I(N__25993));
    LocalMux I__3912 (
            .O(N__25996),
            .I(N__25990));
    LocalMux I__3911 (
            .O(N__25993),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__3910 (
            .O(N__25990),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__3909 (
            .O(N__25985),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__3908 (
            .O(N__25982),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__3907 (
            .O(N__25979),
            .I(N__25975));
    InMux I__3906 (
            .O(N__25978),
            .I(N__25971));
    LocalMux I__3905 (
            .O(N__25975),
            .I(N__25968));
    InMux I__3904 (
            .O(N__25974),
            .I(N__25965));
    LocalMux I__3903 (
            .O(N__25971),
            .I(N__25960));
    Span4Mux_v I__3902 (
            .O(N__25968),
            .I(N__25960));
    LocalMux I__3901 (
            .O(N__25965),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__3900 (
            .O(N__25960),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    InMux I__3899 (
            .O(N__25955),
            .I(N__25952));
    LocalMux I__3898 (
            .O(N__25952),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    CascadeMux I__3897 (
            .O(N__25949),
            .I(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ));
    InMux I__3896 (
            .O(N__25946),
            .I(N__25943));
    LocalMux I__3895 (
            .O(N__25943),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__3894 (
            .O(N__25940),
            .I(N__25936));
    InMux I__3893 (
            .O(N__25939),
            .I(N__25933));
    LocalMux I__3892 (
            .O(N__25936),
            .I(N__25930));
    LocalMux I__3891 (
            .O(N__25933),
            .I(N__25925));
    Span4Mux_h I__3890 (
            .O(N__25930),
            .I(N__25925));
    Odrv4 I__3889 (
            .O(N__25925),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__3888 (
            .O(N__25922),
            .I(N__25918));
    CascadeMux I__3887 (
            .O(N__25921),
            .I(N__25915));
    LocalMux I__3886 (
            .O(N__25918),
            .I(N__25912));
    InMux I__3885 (
            .O(N__25915),
            .I(N__25909));
    Span4Mux_v I__3884 (
            .O(N__25912),
            .I(N__25905));
    LocalMux I__3883 (
            .O(N__25909),
            .I(N__25902));
    InMux I__3882 (
            .O(N__25908),
            .I(N__25899));
    Odrv4 I__3881 (
            .O(N__25905),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__3880 (
            .O(N__25902),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__3879 (
            .O(N__25899),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__3878 (
            .O(N__25892),
            .I(bfn_10_17_0_));
    InMux I__3877 (
            .O(N__25889),
            .I(N__25886));
    LocalMux I__3876 (
            .O(N__25886),
            .I(N__25883));
    Span4Mux_v I__3875 (
            .O(N__25883),
            .I(N__25879));
    InMux I__3874 (
            .O(N__25882),
            .I(N__25876));
    Span4Mux_h I__3873 (
            .O(N__25879),
            .I(N__25872));
    LocalMux I__3872 (
            .O(N__25876),
            .I(N__25869));
    InMux I__3871 (
            .O(N__25875),
            .I(N__25866));
    Odrv4 I__3870 (
            .O(N__25872),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__3869 (
            .O(N__25869),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__3868 (
            .O(N__25866),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__3867 (
            .O(N__25859),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__3866 (
            .O(N__25856),
            .I(N__25849));
    InMux I__3865 (
            .O(N__25855),
            .I(N__25849));
    InMux I__3864 (
            .O(N__25854),
            .I(N__25846));
    LocalMux I__3863 (
            .O(N__25849),
            .I(N__25843));
    LocalMux I__3862 (
            .O(N__25846),
            .I(N__25838));
    Span4Mux_v I__3861 (
            .O(N__25843),
            .I(N__25838));
    Odrv4 I__3860 (
            .O(N__25838),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__3859 (
            .O(N__25835),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__3858 (
            .O(N__25832),
            .I(N__25829));
    InMux I__3857 (
            .O(N__25829),
            .I(N__25825));
    InMux I__3856 (
            .O(N__25828),
            .I(N__25821));
    LocalMux I__3855 (
            .O(N__25825),
            .I(N__25818));
    InMux I__3854 (
            .O(N__25824),
            .I(N__25815));
    LocalMux I__3853 (
            .O(N__25821),
            .I(N__25812));
    Span4Mux_v I__3852 (
            .O(N__25818),
            .I(N__25809));
    LocalMux I__3851 (
            .O(N__25815),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__3850 (
            .O(N__25812),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__3849 (
            .O(N__25809),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__3848 (
            .O(N__25802),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__3847 (
            .O(N__25799),
            .I(N__25796));
    InMux I__3846 (
            .O(N__25796),
            .I(N__25793));
    LocalMux I__3845 (
            .O(N__25793),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__3844 (
            .O(N__25790),
            .I(N__25787));
    LocalMux I__3843 (
            .O(N__25787),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    InMux I__3842 (
            .O(N__25784),
            .I(N__25781));
    LocalMux I__3841 (
            .O(N__25781),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    CascadeMux I__3840 (
            .O(N__25778),
            .I(N__25775));
    InMux I__3839 (
            .O(N__25775),
            .I(N__25772));
    LocalMux I__3838 (
            .O(N__25772),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    InMux I__3837 (
            .O(N__25769),
            .I(N__25766));
    LocalMux I__3836 (
            .O(N__25766),
            .I(N__25763));
    Odrv12 I__3835 (
            .O(N__25763),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    CascadeMux I__3834 (
            .O(N__25760),
            .I(N__25757));
    InMux I__3833 (
            .O(N__25757),
            .I(N__25754));
    LocalMux I__3832 (
            .O(N__25754),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    InMux I__3831 (
            .O(N__25751),
            .I(bfn_10_13_0_));
    CascadeMux I__3830 (
            .O(N__25748),
            .I(N__25745));
    InMux I__3829 (
            .O(N__25745),
            .I(N__25742));
    LocalMux I__3828 (
            .O(N__25742),
            .I(N__25739));
    Span4Mux_h I__3827 (
            .O(N__25739),
            .I(N__25736));
    Span4Mux_h I__3826 (
            .O(N__25736),
            .I(N__25733));
    Odrv4 I__3825 (
            .O(N__25733),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    InMux I__3824 (
            .O(N__25730),
            .I(N__25727));
    LocalMux I__3823 (
            .O(N__25727),
            .I(N__25724));
    Odrv4 I__3822 (
            .O(N__25724),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__3821 (
            .O(N__25721),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    CascadeMux I__3820 (
            .O(N__25718),
            .I(N__25715));
    InMux I__3819 (
            .O(N__25715),
            .I(N__25712));
    LocalMux I__3818 (
            .O(N__25712),
            .I(N__25709));
    Span4Mux_v I__3817 (
            .O(N__25709),
            .I(N__25706));
    Odrv4 I__3816 (
            .O(N__25706),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    InMux I__3815 (
            .O(N__25703),
            .I(N__25700));
    LocalMux I__3814 (
            .O(N__25700),
            .I(N__25697));
    Span4Mux_h I__3813 (
            .O(N__25697),
            .I(N__25694));
    Odrv4 I__3812 (
            .O(N__25694),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__3811 (
            .O(N__25691),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    CascadeMux I__3810 (
            .O(N__25688),
            .I(N__25685));
    InMux I__3809 (
            .O(N__25685),
            .I(N__25682));
    LocalMux I__3808 (
            .O(N__25682),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    InMux I__3807 (
            .O(N__25679),
            .I(N__25676));
    LocalMux I__3806 (
            .O(N__25676),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__3805 (
            .O(N__25673),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    CascadeMux I__3804 (
            .O(N__25670),
            .I(N__25667));
    InMux I__3803 (
            .O(N__25667),
            .I(N__25664));
    LocalMux I__3802 (
            .O(N__25664),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    InMux I__3801 (
            .O(N__25661),
            .I(N__25658));
    LocalMux I__3800 (
            .O(N__25658),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__3799 (
            .O(N__25655),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__3798 (
            .O(N__25652),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    InMux I__3797 (
            .O(N__25649),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    InMux I__3796 (
            .O(N__25646),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__3795 (
            .O(N__25643),
            .I(bfn_10_14_0_));
    CascadeMux I__3794 (
            .O(N__25640),
            .I(N__25637));
    InMux I__3793 (
            .O(N__25637),
            .I(N__25634));
    LocalMux I__3792 (
            .O(N__25634),
            .I(N__25631));
    Odrv4 I__3791 (
            .O(N__25631),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3790 (
            .O(N__25628),
            .I(bfn_10_12_0_));
    CascadeMux I__3789 (
            .O(N__25625),
            .I(N__25622));
    InMux I__3788 (
            .O(N__25622),
            .I(N__25619));
    LocalMux I__3787 (
            .O(N__25619),
            .I(N__25616));
    Span4Mux_h I__3786 (
            .O(N__25616),
            .I(N__25613));
    Span4Mux_h I__3785 (
            .O(N__25613),
            .I(N__25610));
    Odrv4 I__3784 (
            .O(N__25610),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    InMux I__3783 (
            .O(N__25607),
            .I(N__25604));
    LocalMux I__3782 (
            .O(N__25604),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3781 (
            .O(N__25601),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    CascadeMux I__3780 (
            .O(N__25598),
            .I(N__25595));
    InMux I__3779 (
            .O(N__25595),
            .I(N__25592));
    LocalMux I__3778 (
            .O(N__25592),
            .I(N__25589));
    Span4Mux_h I__3777 (
            .O(N__25589),
            .I(N__25586));
    Span4Mux_h I__3776 (
            .O(N__25586),
            .I(N__25583));
    Odrv4 I__3775 (
            .O(N__25583),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    CascadeMux I__3774 (
            .O(N__25580),
            .I(N__25577));
    InMux I__3773 (
            .O(N__25577),
            .I(N__25574));
    LocalMux I__3772 (
            .O(N__25574),
            .I(N__25571));
    Odrv4 I__3771 (
            .O(N__25571),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3770 (
            .O(N__25568),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    CascadeMux I__3769 (
            .O(N__25565),
            .I(N__25562));
    InMux I__3768 (
            .O(N__25562),
            .I(N__25559));
    LocalMux I__3767 (
            .O(N__25559),
            .I(N__25556));
    Span4Mux_v I__3766 (
            .O(N__25556),
            .I(N__25553));
    Odrv4 I__3765 (
            .O(N__25553),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    InMux I__3764 (
            .O(N__25550),
            .I(N__25547));
    LocalMux I__3763 (
            .O(N__25547),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3762 (
            .O(N__25544),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    CascadeMux I__3761 (
            .O(N__25541),
            .I(N__25538));
    InMux I__3760 (
            .O(N__25538),
            .I(N__25535));
    LocalMux I__3759 (
            .O(N__25535),
            .I(N__25532));
    Span4Mux_h I__3758 (
            .O(N__25532),
            .I(N__25529));
    Odrv4 I__3757 (
            .O(N__25529),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    CascadeMux I__3756 (
            .O(N__25526),
            .I(N__25523));
    InMux I__3755 (
            .O(N__25523),
            .I(N__25520));
    LocalMux I__3754 (
            .O(N__25520),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__3753 (
            .O(N__25517),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    CascadeMux I__3752 (
            .O(N__25514),
            .I(N__25511));
    InMux I__3751 (
            .O(N__25511),
            .I(N__25508));
    LocalMux I__3750 (
            .O(N__25508),
            .I(N__25505));
    Odrv4 I__3749 (
            .O(N__25505),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__3748 (
            .O(N__25502),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    InMux I__3747 (
            .O(N__25499),
            .I(N__25496));
    LocalMux I__3746 (
            .O(N__25496),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3745 (
            .O(N__25493),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    CascadeMux I__3744 (
            .O(N__25490),
            .I(N__25487));
    InMux I__3743 (
            .O(N__25487),
            .I(N__25484));
    LocalMux I__3742 (
            .O(N__25484),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3741 (
            .O(N__25481),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    InMux I__3740 (
            .O(N__25478),
            .I(N__25475));
    LocalMux I__3739 (
            .O(N__25475),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3738 (
            .O(N__25472),
            .I(N__25469));
    LocalMux I__3737 (
            .O(N__25469),
            .I(N__25466));
    Odrv4 I__3736 (
            .O(N__25466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ));
    CascadeMux I__3735 (
            .O(N__25463),
            .I(N__25460));
    InMux I__3734 (
            .O(N__25460),
            .I(N__25457));
    LocalMux I__3733 (
            .O(N__25457),
            .I(N__25454));
    Span4Mux_v I__3732 (
            .O(N__25454),
            .I(N__25451));
    Odrv4 I__3731 (
            .O(N__25451),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    InMux I__3730 (
            .O(N__25448),
            .I(N__25445));
    LocalMux I__3729 (
            .O(N__25445),
            .I(N__25442));
    Span4Mux_h I__3728 (
            .O(N__25442),
            .I(N__25439));
    Odrv4 I__3727 (
            .O(N__25439),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3726 (
            .O(N__25436),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__3725 (
            .O(N__25433),
            .I(N__25430));
    LocalMux I__3724 (
            .O(N__25430),
            .I(N__25427));
    Odrv4 I__3723 (
            .O(N__25427),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ));
    CascadeMux I__3722 (
            .O(N__25424),
            .I(N__25421));
    InMux I__3721 (
            .O(N__25421),
            .I(N__25418));
    LocalMux I__3720 (
            .O(N__25418),
            .I(N__25415));
    Span4Mux_v I__3719 (
            .O(N__25415),
            .I(N__25412));
    Odrv4 I__3718 (
            .O(N__25412),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    InMux I__3717 (
            .O(N__25409),
            .I(N__25406));
    LocalMux I__3716 (
            .O(N__25406),
            .I(N__25403));
    Span4Mux_h I__3715 (
            .O(N__25403),
            .I(N__25400));
    Odrv4 I__3714 (
            .O(N__25400),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__3713 (
            .O(N__25397),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    InMux I__3712 (
            .O(N__25394),
            .I(N__25391));
    LocalMux I__3711 (
            .O(N__25391),
            .I(N__25388));
    Odrv4 I__3710 (
            .O(N__25388),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ));
    CascadeMux I__3709 (
            .O(N__25385),
            .I(N__25382));
    InMux I__3708 (
            .O(N__25382),
            .I(N__25379));
    LocalMux I__3707 (
            .O(N__25379),
            .I(N__25376));
    Span4Mux_v I__3706 (
            .O(N__25376),
            .I(N__25373));
    Odrv4 I__3705 (
            .O(N__25373),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    InMux I__3704 (
            .O(N__25370),
            .I(N__25367));
    LocalMux I__3703 (
            .O(N__25367),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__3702 (
            .O(N__25364),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__3701 (
            .O(N__25361),
            .I(N__25358));
    LocalMux I__3700 (
            .O(N__25358),
            .I(N__25355));
    Odrv4 I__3699 (
            .O(N__25355),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ));
    InMux I__3698 (
            .O(N__25352),
            .I(N__25349));
    LocalMux I__3697 (
            .O(N__25349),
            .I(N__25346));
    Odrv4 I__3696 (
            .O(N__25346),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3695 (
            .O(N__25343),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    CascadeMux I__3694 (
            .O(N__25340),
            .I(N__25337));
    InMux I__3693 (
            .O(N__25337),
            .I(N__25334));
    LocalMux I__3692 (
            .O(N__25334),
            .I(N__25331));
    Span4Mux_h I__3691 (
            .O(N__25331),
            .I(N__25328));
    Odrv4 I__3690 (
            .O(N__25328),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    InMux I__3689 (
            .O(N__25325),
            .I(N__25322));
    LocalMux I__3688 (
            .O(N__25322),
            .I(N__25319));
    Span4Mux_h I__3687 (
            .O(N__25319),
            .I(N__25316));
    Odrv4 I__3686 (
            .O(N__25316),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3685 (
            .O(N__25313),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    CascadeMux I__3684 (
            .O(N__25310),
            .I(N__25307));
    InMux I__3683 (
            .O(N__25307),
            .I(N__25304));
    LocalMux I__3682 (
            .O(N__25304),
            .I(N__25301));
    Span4Mux_v I__3681 (
            .O(N__25301),
            .I(N__25298));
    Odrv4 I__3680 (
            .O(N__25298),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    CascadeMux I__3679 (
            .O(N__25295),
            .I(N__25292));
    InMux I__3678 (
            .O(N__25292),
            .I(N__25289));
    LocalMux I__3677 (
            .O(N__25289),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3676 (
            .O(N__25286),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    InMux I__3675 (
            .O(N__25283),
            .I(N__25280));
    LocalMux I__3674 (
            .O(N__25280),
            .I(N__25277));
    Odrv4 I__3673 (
            .O(N__25277),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__3672 (
            .O(N__25274),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    CascadeMux I__3671 (
            .O(N__25271),
            .I(N__25268));
    InMux I__3670 (
            .O(N__25268),
            .I(N__25265));
    LocalMux I__3669 (
            .O(N__25265),
            .I(N__25262));
    Span4Mux_h I__3668 (
            .O(N__25262),
            .I(N__25259));
    Odrv4 I__3667 (
            .O(N__25259),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    CascadeMux I__3666 (
            .O(N__25256),
            .I(N__25253));
    InMux I__3665 (
            .O(N__25253),
            .I(N__25249));
    InMux I__3664 (
            .O(N__25252),
            .I(N__25246));
    LocalMux I__3663 (
            .O(N__25249),
            .I(N__25241));
    LocalMux I__3662 (
            .O(N__25246),
            .I(N__25241));
    Odrv4 I__3661 (
            .O(N__25241),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__3660 (
            .O(N__25238),
            .I(N__25235));
    InMux I__3659 (
            .O(N__25235),
            .I(N__25232));
    LocalMux I__3658 (
            .O(N__25232),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ));
    InMux I__3657 (
            .O(N__25229),
            .I(N__25226));
    LocalMux I__3656 (
            .O(N__25226),
            .I(N__25223));
    Odrv4 I__3655 (
            .O(N__25223),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ));
    InMux I__3654 (
            .O(N__25220),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__3653 (
            .O(N__25217),
            .I(N__25214));
    LocalMux I__3652 (
            .O(N__25214),
            .I(N__25211));
    Odrv4 I__3651 (
            .O(N__25211),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ));
    CascadeMux I__3650 (
            .O(N__25208),
            .I(N__25205));
    InMux I__3649 (
            .O(N__25205),
            .I(N__25202));
    LocalMux I__3648 (
            .O(N__25202),
            .I(N__25199));
    Odrv4 I__3647 (
            .O(N__25199),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    InMux I__3646 (
            .O(N__25196),
            .I(N__25193));
    LocalMux I__3645 (
            .O(N__25193),
            .I(N__25190));
    Span4Mux_v I__3644 (
            .O(N__25190),
            .I(N__25187));
    Odrv4 I__3643 (
            .O(N__25187),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__3642 (
            .O(N__25184),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__3641 (
            .O(N__25181),
            .I(N__25178));
    LocalMux I__3640 (
            .O(N__25178),
            .I(N__25175));
    Odrv4 I__3639 (
            .O(N__25175),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ));
    CascadeMux I__3638 (
            .O(N__25172),
            .I(N__25169));
    InMux I__3637 (
            .O(N__25169),
            .I(N__25166));
    LocalMux I__3636 (
            .O(N__25166),
            .I(N__25163));
    Odrv4 I__3635 (
            .O(N__25163),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    InMux I__3634 (
            .O(N__25160),
            .I(N__25157));
    LocalMux I__3633 (
            .O(N__25157),
            .I(N__25154));
    Odrv4 I__3632 (
            .O(N__25154),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__3631 (
            .O(N__25151),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__3630 (
            .O(N__25148),
            .I(N__25145));
    LocalMux I__3629 (
            .O(N__25145),
            .I(N__25142));
    Odrv4 I__3628 (
            .O(N__25142),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ));
    CascadeMux I__3627 (
            .O(N__25139),
            .I(N__25136));
    InMux I__3626 (
            .O(N__25136),
            .I(N__25133));
    LocalMux I__3625 (
            .O(N__25133),
            .I(N__25130));
    Odrv4 I__3624 (
            .O(N__25130),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    InMux I__3623 (
            .O(N__25127),
            .I(N__25124));
    LocalMux I__3622 (
            .O(N__25124),
            .I(N__25121));
    Odrv4 I__3621 (
            .O(N__25121),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__3620 (
            .O(N__25118),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__3619 (
            .O(N__25115),
            .I(N__25112));
    LocalMux I__3618 (
            .O(N__25112),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ));
    CascadeMux I__3617 (
            .O(N__25109),
            .I(N__25106));
    InMux I__3616 (
            .O(N__25106),
            .I(N__25103));
    LocalMux I__3615 (
            .O(N__25103),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    InMux I__3614 (
            .O(N__25100),
            .I(N__25097));
    LocalMux I__3613 (
            .O(N__25097),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__3612 (
            .O(N__25094),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__3611 (
            .O(N__25091),
            .I(N__25088));
    LocalMux I__3610 (
            .O(N__25088),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ));
    CascadeMux I__3609 (
            .O(N__25085),
            .I(N__25082));
    InMux I__3608 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__3607 (
            .O(N__25079),
            .I(N__25076));
    Span4Mux_h I__3606 (
            .O(N__25076),
            .I(N__25073));
    Odrv4 I__3605 (
            .O(N__25073),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    InMux I__3604 (
            .O(N__25070),
            .I(N__25067));
    LocalMux I__3603 (
            .O(N__25067),
            .I(N__25064));
    Odrv4 I__3602 (
            .O(N__25064),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__3601 (
            .O(N__25061),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__3600 (
            .O(N__25058),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__3599 (
            .O(N__25055),
            .I(N__25052));
    LocalMux I__3598 (
            .O(N__25052),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ));
    CascadeMux I__3597 (
            .O(N__25049),
            .I(N__25046));
    InMux I__3596 (
            .O(N__25046),
            .I(N__25043));
    LocalMux I__3595 (
            .O(N__25043),
            .I(N__25040));
    Odrv4 I__3594 (
            .O(N__25040),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    InMux I__3593 (
            .O(N__25037),
            .I(N__25034));
    LocalMux I__3592 (
            .O(N__25034),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__3591 (
            .O(N__25031),
            .I(bfn_10_11_0_));
    CascadeMux I__3590 (
            .O(N__25028),
            .I(N__25025));
    InMux I__3589 (
            .O(N__25025),
            .I(N__25021));
    InMux I__3588 (
            .O(N__25024),
            .I(N__25018));
    LocalMux I__3587 (
            .O(N__25021),
            .I(N__25013));
    LocalMux I__3586 (
            .O(N__25018),
            .I(N__25010));
    InMux I__3585 (
            .O(N__25017),
            .I(N__25006));
    InMux I__3584 (
            .O(N__25016),
            .I(N__25003));
    Span4Mux_h I__3583 (
            .O(N__25013),
            .I(N__25000));
    Span4Mux_v I__3582 (
            .O(N__25010),
            .I(N__24997));
    InMux I__3581 (
            .O(N__25009),
            .I(N__24994));
    LocalMux I__3580 (
            .O(N__25006),
            .I(N__24989));
    LocalMux I__3579 (
            .O(N__25003),
            .I(N__24989));
    Odrv4 I__3578 (
            .O(N__25000),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__3577 (
            .O(N__24997),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__3576 (
            .O(N__24994),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__3575 (
            .O(N__24989),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__3574 (
            .O(N__24980),
            .I(N__24977));
    InMux I__3573 (
            .O(N__24977),
            .I(N__24973));
    InMux I__3572 (
            .O(N__24976),
            .I(N__24970));
    LocalMux I__3571 (
            .O(N__24973),
            .I(N__24966));
    LocalMux I__3570 (
            .O(N__24970),
            .I(N__24961));
    InMux I__3569 (
            .O(N__24969),
            .I(N__24958));
    Span4Mux_h I__3568 (
            .O(N__24966),
            .I(N__24955));
    InMux I__3567 (
            .O(N__24965),
            .I(N__24952));
    InMux I__3566 (
            .O(N__24964),
            .I(N__24949));
    Span4Mux_v I__3565 (
            .O(N__24961),
            .I(N__24944));
    LocalMux I__3564 (
            .O(N__24958),
            .I(N__24944));
    Odrv4 I__3563 (
            .O(N__24955),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3562 (
            .O(N__24952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3561 (
            .O(N__24949),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__3560 (
            .O(N__24944),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__3559 (
            .O(N__24935),
            .I(N__24930));
    InMux I__3558 (
            .O(N__24934),
            .I(N__24927));
    CascadeMux I__3557 (
            .O(N__24933),
            .I(N__24922));
    LocalMux I__3556 (
            .O(N__24930),
            .I(N__24919));
    LocalMux I__3555 (
            .O(N__24927),
            .I(N__24916));
    InMux I__3554 (
            .O(N__24926),
            .I(N__24911));
    InMux I__3553 (
            .O(N__24925),
            .I(N__24911));
    InMux I__3552 (
            .O(N__24922),
            .I(N__24908));
    Span4Mux_h I__3551 (
            .O(N__24919),
            .I(N__24905));
    Span4Mux_h I__3550 (
            .O(N__24916),
            .I(N__24900));
    LocalMux I__3549 (
            .O(N__24911),
            .I(N__24900));
    LocalMux I__3548 (
            .O(N__24908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3547 (
            .O(N__24905),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3546 (
            .O(N__24900),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__3545 (
            .O(N__24893),
            .I(N__24890));
    InMux I__3544 (
            .O(N__24890),
            .I(N__24887));
    LocalMux I__3543 (
            .O(N__24887),
            .I(N__24881));
    InMux I__3542 (
            .O(N__24886),
            .I(N__24877));
    InMux I__3541 (
            .O(N__24885),
            .I(N__24874));
    CascadeMux I__3540 (
            .O(N__24884),
            .I(N__24871));
    Span4Mux_v I__3539 (
            .O(N__24881),
            .I(N__24868));
    InMux I__3538 (
            .O(N__24880),
            .I(N__24865));
    LocalMux I__3537 (
            .O(N__24877),
            .I(N__24860));
    LocalMux I__3536 (
            .O(N__24874),
            .I(N__24860));
    InMux I__3535 (
            .O(N__24871),
            .I(N__24857));
    Odrv4 I__3534 (
            .O(N__24868),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3533 (
            .O(N__24865),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__3532 (
            .O(N__24860),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3531 (
            .O(N__24857),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__3530 (
            .O(N__24848),
            .I(N__24845));
    InMux I__3529 (
            .O(N__24845),
            .I(N__24841));
    InMux I__3528 (
            .O(N__24844),
            .I(N__24838));
    LocalMux I__3527 (
            .O(N__24841),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_16 ));
    LocalMux I__3526 (
            .O(N__24838),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_16 ));
    InMux I__3525 (
            .O(N__24833),
            .I(N__24828));
    InMux I__3524 (
            .O(N__24832),
            .I(N__24825));
    InMux I__3523 (
            .O(N__24831),
            .I(N__24822));
    LocalMux I__3522 (
            .O(N__24828),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__3521 (
            .O(N__24825),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__3520 (
            .O(N__24822),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__3519 (
            .O(N__24815),
            .I(N__24810));
    InMux I__3518 (
            .O(N__24814),
            .I(N__24807));
    InMux I__3517 (
            .O(N__24813),
            .I(N__24804));
    LocalMux I__3516 (
            .O(N__24810),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__3515 (
            .O(N__24807),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__3514 (
            .O(N__24804),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    CascadeMux I__3513 (
            .O(N__24797),
            .I(N__24794));
    InMux I__3512 (
            .O(N__24794),
            .I(N__24791));
    LocalMux I__3511 (
            .O(N__24791),
            .I(N__24788));
    Span4Mux_v I__3510 (
            .O(N__24788),
            .I(N__24785));
    Odrv4 I__3509 (
            .O(N__24785),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__3508 (
            .O(N__24782),
            .I(N__24779));
    LocalMux I__3507 (
            .O(N__24779),
            .I(N__24775));
    InMux I__3506 (
            .O(N__24778),
            .I(N__24772));
    Span4Mux_v I__3505 (
            .O(N__24775),
            .I(N__24768));
    LocalMux I__3504 (
            .O(N__24772),
            .I(N__24765));
    CascadeMux I__3503 (
            .O(N__24771),
            .I(N__24762));
    Span4Mux_h I__3502 (
            .O(N__24768),
            .I(N__24756));
    Span4Mux_v I__3501 (
            .O(N__24765),
            .I(N__24756));
    InMux I__3500 (
            .O(N__24762),
            .I(N__24751));
    InMux I__3499 (
            .O(N__24761),
            .I(N__24751));
    Odrv4 I__3498 (
            .O(N__24756),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__3497 (
            .O(N__24751),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__3496 (
            .O(N__24746),
            .I(N__24741));
    InMux I__3495 (
            .O(N__24745),
            .I(N__24738));
    CascadeMux I__3494 (
            .O(N__24744),
            .I(N__24735));
    LocalMux I__3493 (
            .O(N__24741),
            .I(N__24732));
    LocalMux I__3492 (
            .O(N__24738),
            .I(N__24729));
    InMux I__3491 (
            .O(N__24735),
            .I(N__24724));
    Span12Mux_v I__3490 (
            .O(N__24732),
            .I(N__24721));
    Span4Mux_v I__3489 (
            .O(N__24729),
            .I(N__24718));
    InMux I__3488 (
            .O(N__24728),
            .I(N__24715));
    InMux I__3487 (
            .O(N__24727),
            .I(N__24712));
    LocalMux I__3486 (
            .O(N__24724),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__3485 (
            .O(N__24721),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3484 (
            .O(N__24718),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__3483 (
            .O(N__24715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__3482 (
            .O(N__24712),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__3481 (
            .O(N__24701),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9_cascade_ ));
    InMux I__3480 (
            .O(N__24698),
            .I(N__24695));
    LocalMux I__3479 (
            .O(N__24695),
            .I(N__24692));
    Odrv4 I__3478 (
            .O(N__24692),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ));
    InMux I__3477 (
            .O(N__24689),
            .I(N__24683));
    InMux I__3476 (
            .O(N__24688),
            .I(N__24683));
    LocalMux I__3475 (
            .O(N__24683),
            .I(\delay_measurement_inst.elapsed_time_hc_28 ));
    InMux I__3474 (
            .O(N__24680),
            .I(N__24677));
    LocalMux I__3473 (
            .O(N__24677),
            .I(\delay_measurement_inst.N_52 ));
    InMux I__3472 (
            .O(N__24674),
            .I(N__24671));
    LocalMux I__3471 (
            .O(N__24671),
            .I(N__24668));
    Glb2LocalMux I__3470 (
            .O(N__24668),
            .I(N__24665));
    GlobalMux I__3469 (
            .O(N__24665),
            .I(clk_12mhz));
    IoInMux I__3468 (
            .O(N__24662),
            .I(N__24659));
    LocalMux I__3467 (
            .O(N__24659),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__3466 (
            .O(N__24656),
            .I(N__24653));
    LocalMux I__3465 (
            .O(N__24653),
            .I(N__24650));
    Span4Mux_h I__3464 (
            .O(N__24650),
            .I(N__24647));
    Odrv4 I__3463 (
            .O(N__24647),
            .I(il_min_comp1_c));
    InMux I__3462 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__3461 (
            .O(N__24641),
            .I(N__24638));
    Span4Mux_h I__3460 (
            .O(N__24638),
            .I(N__24635));
    Odrv4 I__3459 (
            .O(N__24635),
            .I(il_max_comp1_D1));
    InMux I__3458 (
            .O(N__24632),
            .I(N__24629));
    LocalMux I__3457 (
            .O(N__24629),
            .I(il_min_comp1_D1));
    InMux I__3456 (
            .O(N__24626),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__3455 (
            .O(N__24623),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__3454 (
            .O(N__24620),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__3453 (
            .O(N__24617),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__3452 (
            .O(N__24614),
            .I(bfn_9_22_0_));
    InMux I__3451 (
            .O(N__24611),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__3450 (
            .O(N__24608),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__3449 (
            .O(N__24605),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__3448 (
            .O(N__24602),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__3447 (
            .O(N__24599),
            .I(N__24584));
    CEMux I__3446 (
            .O(N__24598),
            .I(N__24584));
    CEMux I__3445 (
            .O(N__24597),
            .I(N__24584));
    CEMux I__3444 (
            .O(N__24596),
            .I(N__24584));
    CEMux I__3443 (
            .O(N__24595),
            .I(N__24584));
    GlobalMux I__3442 (
            .O(N__24584),
            .I(N__24581));
    gio2CtrlBuf I__3441 (
            .O(N__24581),
            .I(\delay_measurement_inst.delay_hc_timer.N_302_i_g ));
    InMux I__3440 (
            .O(N__24578),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__3439 (
            .O(N__24575),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__3438 (
            .O(N__24572),
            .I(N__24567));
    InMux I__3437 (
            .O(N__24571),
            .I(N__24564));
    InMux I__3436 (
            .O(N__24570),
            .I(N__24559));
    InMux I__3435 (
            .O(N__24567),
            .I(N__24559));
    LocalMux I__3434 (
            .O(N__24564),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__3433 (
            .O(N__24559),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__3432 (
            .O(N__24554),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__3431 (
            .O(N__24551),
            .I(N__24547));
    InMux I__3430 (
            .O(N__24550),
            .I(N__24543));
    LocalMux I__3429 (
            .O(N__24547),
            .I(N__24540));
    InMux I__3428 (
            .O(N__24546),
            .I(N__24537));
    LocalMux I__3427 (
            .O(N__24543),
            .I(N__24534));
    Odrv4 I__3426 (
            .O(N__24540),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__3425 (
            .O(N__24537),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    Odrv4 I__3424 (
            .O(N__24534),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__3423 (
            .O(N__24527),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__3422 (
            .O(N__24524),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__3421 (
            .O(N__24521),
            .I(N__24517));
    InMux I__3420 (
            .O(N__24520),
            .I(N__24513));
    InMux I__3419 (
            .O(N__24517),
            .I(N__24510));
    InMux I__3418 (
            .O(N__24516),
            .I(N__24507));
    LocalMux I__3417 (
            .O(N__24513),
            .I(N__24502));
    LocalMux I__3416 (
            .O(N__24510),
            .I(N__24502));
    LocalMux I__3415 (
            .O(N__24507),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__3414 (
            .O(N__24502),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__3413 (
            .O(N__24497),
            .I(bfn_9_21_0_));
    InMux I__3412 (
            .O(N__24494),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__3411 (
            .O(N__24491),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__3410 (
            .O(N__24488),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__3409 (
            .O(N__24485),
            .I(N__24481));
    InMux I__3408 (
            .O(N__24484),
            .I(N__24478));
    LocalMux I__3407 (
            .O(N__24481),
            .I(N__24473));
    LocalMux I__3406 (
            .O(N__24478),
            .I(N__24473));
    Span4Mux_v I__3405 (
            .O(N__24473),
            .I(N__24468));
    InMux I__3404 (
            .O(N__24472),
            .I(N__24463));
    InMux I__3403 (
            .O(N__24471),
            .I(N__24463));
    Odrv4 I__3402 (
            .O(N__24468),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__3401 (
            .O(N__24463),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__3400 (
            .O(N__24458),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__3399 (
            .O(N__24455),
            .I(N__24452));
    LocalMux I__3398 (
            .O(N__24452),
            .I(N__24446));
    InMux I__3397 (
            .O(N__24451),
            .I(N__24443));
    InMux I__3396 (
            .O(N__24450),
            .I(N__24438));
    InMux I__3395 (
            .O(N__24449),
            .I(N__24438));
    Odrv4 I__3394 (
            .O(N__24446),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__3393 (
            .O(N__24443),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__3392 (
            .O(N__24438),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__3391 (
            .O(N__24431),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__3390 (
            .O(N__24428),
            .I(N__24424));
    InMux I__3389 (
            .O(N__24427),
            .I(N__24421));
    LocalMux I__3388 (
            .O(N__24424),
            .I(N__24416));
    LocalMux I__3387 (
            .O(N__24421),
            .I(N__24416));
    Span4Mux_h I__3386 (
            .O(N__24416),
            .I(N__24411));
    InMux I__3385 (
            .O(N__24415),
            .I(N__24408));
    InMux I__3384 (
            .O(N__24414),
            .I(N__24405));
    Odrv4 I__3383 (
            .O(N__24411),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__3382 (
            .O(N__24408),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__3381 (
            .O(N__24405),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__3380 (
            .O(N__24398),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__3379 (
            .O(N__24395),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__3378 (
            .O(N__24392),
            .I(N__24386));
    InMux I__3377 (
            .O(N__24391),
            .I(N__24386));
    LocalMux I__3376 (
            .O(N__24386),
            .I(N__24382));
    InMux I__3375 (
            .O(N__24385),
            .I(N__24379));
    Span4Mux_h I__3374 (
            .O(N__24382),
            .I(N__24376));
    LocalMux I__3373 (
            .O(N__24379),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    Odrv4 I__3372 (
            .O(N__24376),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__3371 (
            .O(N__24371),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__3370 (
            .O(N__24368),
            .I(N__24365));
    LocalMux I__3369 (
            .O(N__24365),
            .I(N__24362));
    Span4Mux_h I__3368 (
            .O(N__24362),
            .I(N__24357));
    InMux I__3367 (
            .O(N__24361),
            .I(N__24354));
    InMux I__3366 (
            .O(N__24360),
            .I(N__24351));
    Odrv4 I__3365 (
            .O(N__24357),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    LocalMux I__3364 (
            .O(N__24354),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    LocalMux I__3363 (
            .O(N__24351),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__3362 (
            .O(N__24344),
            .I(bfn_9_20_0_));
    InMux I__3361 (
            .O(N__24341),
            .I(N__24338));
    LocalMux I__3360 (
            .O(N__24338),
            .I(N__24333));
    CascadeMux I__3359 (
            .O(N__24337),
            .I(N__24330));
    CascadeMux I__3358 (
            .O(N__24336),
            .I(N__24327));
    Span4Mux_v I__3357 (
            .O(N__24333),
            .I(N__24324));
    InMux I__3356 (
            .O(N__24330),
            .I(N__24321));
    InMux I__3355 (
            .O(N__24327),
            .I(N__24318));
    Odrv4 I__3354 (
            .O(N__24324),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    LocalMux I__3353 (
            .O(N__24321),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    LocalMux I__3352 (
            .O(N__24318),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__3351 (
            .O(N__24311),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__3350 (
            .O(N__24308),
            .I(N__24305));
    LocalMux I__3349 (
            .O(N__24305),
            .I(N__24300));
    InMux I__3348 (
            .O(N__24304),
            .I(N__24295));
    InMux I__3347 (
            .O(N__24303),
            .I(N__24295));
    Odrv4 I__3346 (
            .O(N__24300),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__3345 (
            .O(N__24295),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__3344 (
            .O(N__24290),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__3343 (
            .O(N__24287),
            .I(N__24281));
    InMux I__3342 (
            .O(N__24286),
            .I(N__24276));
    InMux I__3341 (
            .O(N__24285),
            .I(N__24276));
    InMux I__3340 (
            .O(N__24284),
            .I(N__24273));
    LocalMux I__3339 (
            .O(N__24281),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__3338 (
            .O(N__24276),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__3337 (
            .O(N__24273),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    CascadeMux I__3336 (
            .O(N__24266),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt30_cascade_ ));
    CascadeMux I__3335 (
            .O(N__24263),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1_cascade_ ));
    InMux I__3334 (
            .O(N__24260),
            .I(N__24257));
    LocalMux I__3333 (
            .O(N__24257),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt14_0 ));
    InMux I__3332 (
            .O(N__24254),
            .I(N__24251));
    LocalMux I__3331 (
            .O(N__24251),
            .I(\delay_measurement_inst.N_41 ));
    InMux I__3330 (
            .O(N__24248),
            .I(N__24245));
    LocalMux I__3329 (
            .O(N__24245),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ));
    InMux I__3328 (
            .O(N__24242),
            .I(N__24235));
    InMux I__3327 (
            .O(N__24241),
            .I(N__24235));
    InMux I__3326 (
            .O(N__24240),
            .I(N__24232));
    LocalMux I__3325 (
            .O(N__24235),
            .I(N__24229));
    LocalMux I__3324 (
            .O(N__24232),
            .I(N__24224));
    Span4Mux_h I__3323 (
            .O(N__24229),
            .I(N__24224));
    Odrv4 I__3322 (
            .O(N__24224),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__3321 (
            .O(N__24221),
            .I(N__24216));
    InMux I__3320 (
            .O(N__24220),
            .I(N__24213));
    InMux I__3319 (
            .O(N__24219),
            .I(N__24210));
    LocalMux I__3318 (
            .O(N__24216),
            .I(N__24207));
    LocalMux I__3317 (
            .O(N__24213),
            .I(N__24204));
    LocalMux I__3316 (
            .O(N__24210),
            .I(N__24197));
    Span4Mux_v I__3315 (
            .O(N__24207),
            .I(N__24197));
    Span4Mux_h I__3314 (
            .O(N__24204),
            .I(N__24197));
    Odrv4 I__3313 (
            .O(N__24197),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__3312 (
            .O(N__24194),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__3311 (
            .O(N__24191),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__3310 (
            .O(N__24188),
            .I(N__24184));
    InMux I__3309 (
            .O(N__24187),
            .I(N__24181));
    LocalMux I__3308 (
            .O(N__24184),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3307 (
            .O(N__24181),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__3306 (
            .O(N__24176),
            .I(N__24173));
    LocalMux I__3305 (
            .O(N__24173),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__3304 (
            .O(N__24170),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__3303 (
            .O(N__24167),
            .I(N__24163));
    InMux I__3302 (
            .O(N__24166),
            .I(N__24160));
    LocalMux I__3301 (
            .O(N__24163),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3300 (
            .O(N__24160),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3299 (
            .O(N__24155),
            .I(N__24152));
    LocalMux I__3298 (
            .O(N__24152),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__3297 (
            .O(N__24149),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__3296 (
            .O(N__24146),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__3295 (
            .O(N__24143),
            .I(N__24139));
    InMux I__3294 (
            .O(N__24142),
            .I(N__24136));
    LocalMux I__3293 (
            .O(N__24139),
            .I(N__24133));
    LocalMux I__3292 (
            .O(N__24136),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__3291 (
            .O(N__24133),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__3290 (
            .O(N__24128),
            .I(N__24125));
    LocalMux I__3289 (
            .O(N__24125),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__3288 (
            .O(N__24122),
            .I(bfn_9_16_0_));
    InMux I__3287 (
            .O(N__24119),
            .I(N__24115));
    InMux I__3286 (
            .O(N__24118),
            .I(N__24112));
    LocalMux I__3285 (
            .O(N__24115),
            .I(N__24109));
    LocalMux I__3284 (
            .O(N__24112),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__3283 (
            .O(N__24109),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__3282 (
            .O(N__24104),
            .I(N__24101));
    LocalMux I__3281 (
            .O(N__24101),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__3280 (
            .O(N__24098),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__3279 (
            .O(N__24095),
            .I(N__24091));
    InMux I__3278 (
            .O(N__24094),
            .I(N__24088));
    LocalMux I__3277 (
            .O(N__24091),
            .I(N__24085));
    LocalMux I__3276 (
            .O(N__24088),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__3275 (
            .O(N__24085),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__3274 (
            .O(N__24080),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__3273 (
            .O(N__24077),
            .I(N__24074));
    LocalMux I__3272 (
            .O(N__24074),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    CascadeMux I__3271 (
            .O(N__24071),
            .I(N__24068));
    InMux I__3270 (
            .O(N__24068),
            .I(N__24065));
    LocalMux I__3269 (
            .O(N__24065),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    InMux I__3268 (
            .O(N__24062),
            .I(N__24058));
    InMux I__3267 (
            .O(N__24061),
            .I(N__24055));
    LocalMux I__3266 (
            .O(N__24058),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3265 (
            .O(N__24055),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3264 (
            .O(N__24050),
            .I(N__24047));
    LocalMux I__3263 (
            .O(N__24047),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__3262 (
            .O(N__24044),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__3261 (
            .O(N__24041),
            .I(N__24037));
    InMux I__3260 (
            .O(N__24040),
            .I(N__24034));
    LocalMux I__3259 (
            .O(N__24037),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3258 (
            .O(N__24034),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3257 (
            .O(N__24029),
            .I(N__24026));
    LocalMux I__3256 (
            .O(N__24026),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__3255 (
            .O(N__24023),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__3254 (
            .O(N__24020),
            .I(N__24016));
    InMux I__3253 (
            .O(N__24019),
            .I(N__24013));
    LocalMux I__3252 (
            .O(N__24016),
            .I(N__24010));
    LocalMux I__3251 (
            .O(N__24013),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__3250 (
            .O(N__24010),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3249 (
            .O(N__24005),
            .I(N__24002));
    LocalMux I__3248 (
            .O(N__24002),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__3247 (
            .O(N__23999),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__3246 (
            .O(N__23996),
            .I(N__23992));
    InMux I__3245 (
            .O(N__23995),
            .I(N__23989));
    LocalMux I__3244 (
            .O(N__23992),
            .I(N__23986));
    LocalMux I__3243 (
            .O(N__23989),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__3242 (
            .O(N__23986),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3241 (
            .O(N__23981),
            .I(N__23978));
    LocalMux I__3240 (
            .O(N__23978),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__3239 (
            .O(N__23975),
            .I(bfn_9_15_0_));
    InMux I__3238 (
            .O(N__23972),
            .I(N__23968));
    InMux I__3237 (
            .O(N__23971),
            .I(N__23965));
    LocalMux I__3236 (
            .O(N__23968),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3235 (
            .O(N__23965),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__3234 (
            .O(N__23960),
            .I(N__23957));
    LocalMux I__3233 (
            .O(N__23957),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__3232 (
            .O(N__23954),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__3231 (
            .O(N__23951),
            .I(N__23947));
    InMux I__3230 (
            .O(N__23950),
            .I(N__23944));
    LocalMux I__3229 (
            .O(N__23947),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3228 (
            .O(N__23944),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3227 (
            .O(N__23939),
            .I(N__23936));
    LocalMux I__3226 (
            .O(N__23936),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__3225 (
            .O(N__23933),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__3224 (
            .O(N__23930),
            .I(N__23926));
    InMux I__3223 (
            .O(N__23929),
            .I(N__23923));
    LocalMux I__3222 (
            .O(N__23926),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3221 (
            .O(N__23923),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3220 (
            .O(N__23918),
            .I(N__23915));
    LocalMux I__3219 (
            .O(N__23915),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__3218 (
            .O(N__23912),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__3217 (
            .O(N__23909),
            .I(N__23905));
    InMux I__3216 (
            .O(N__23908),
            .I(N__23902));
    LocalMux I__3215 (
            .O(N__23905),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3214 (
            .O(N__23902),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__3213 (
            .O(N__23897),
            .I(N__23894));
    LocalMux I__3212 (
            .O(N__23894),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__3211 (
            .O(N__23891),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__3210 (
            .O(N__23888),
            .I(N__23885));
    LocalMux I__3209 (
            .O(N__23885),
            .I(N__23882));
    Span4Mux_h I__3208 (
            .O(N__23882),
            .I(N__23879));
    Odrv4 I__3207 (
            .O(N__23879),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    CascadeMux I__3206 (
            .O(N__23876),
            .I(N__23873));
    InMux I__3205 (
            .O(N__23873),
            .I(N__23869));
    InMux I__3204 (
            .O(N__23872),
            .I(N__23865));
    LocalMux I__3203 (
            .O(N__23869),
            .I(N__23862));
    InMux I__3202 (
            .O(N__23868),
            .I(N__23859));
    LocalMux I__3201 (
            .O(N__23865),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3200 (
            .O(N__23862),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__3199 (
            .O(N__23859),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__3198 (
            .O(N__23852),
            .I(N__23848));
    InMux I__3197 (
            .O(N__23851),
            .I(N__23845));
    LocalMux I__3196 (
            .O(N__23848),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3195 (
            .O(N__23845),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__3194 (
            .O(N__23840),
            .I(N__23837));
    LocalMux I__3193 (
            .O(N__23837),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__3192 (
            .O(N__23834),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__3191 (
            .O(N__23831),
            .I(N__23827));
    InMux I__3190 (
            .O(N__23830),
            .I(N__23824));
    LocalMux I__3189 (
            .O(N__23827),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3188 (
            .O(N__23824),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__3187 (
            .O(N__23819),
            .I(N__23816));
    LocalMux I__3186 (
            .O(N__23816),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__3185 (
            .O(N__23813),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    CascadeMux I__3184 (
            .O(N__23810),
            .I(N__23807));
    InMux I__3183 (
            .O(N__23807),
            .I(N__23803));
    InMux I__3182 (
            .O(N__23806),
            .I(N__23800));
    LocalMux I__3181 (
            .O(N__23803),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3180 (
            .O(N__23800),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3179 (
            .O(N__23795),
            .I(N__23792));
    LocalMux I__3178 (
            .O(N__23792),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__3177 (
            .O(N__23789),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__3176 (
            .O(N__23786),
            .I(N__23782));
    InMux I__3175 (
            .O(N__23785),
            .I(N__23779));
    LocalMux I__3174 (
            .O(N__23782),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3173 (
            .O(N__23779),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__3172 (
            .O(N__23774),
            .I(N__23771));
    LocalMux I__3171 (
            .O(N__23771),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__3170 (
            .O(N__23768),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    CascadeMux I__3169 (
            .O(N__23765),
            .I(N__23762));
    InMux I__3168 (
            .O(N__23762),
            .I(N__23759));
    LocalMux I__3167 (
            .O(N__23759),
            .I(N__23756));
    Span4Mux_v I__3166 (
            .O(N__23756),
            .I(N__23753));
    Odrv4 I__3165 (
            .O(N__23753),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__3164 (
            .O(N__23750),
            .I(N__23747));
    LocalMux I__3163 (
            .O(N__23747),
            .I(N__23744));
    Span4Mux_h I__3162 (
            .O(N__23744),
            .I(N__23739));
    InMux I__3161 (
            .O(N__23743),
            .I(N__23736));
    InMux I__3160 (
            .O(N__23742),
            .I(N__23733));
    Span4Mux_h I__3159 (
            .O(N__23739),
            .I(N__23730));
    LocalMux I__3158 (
            .O(N__23736),
            .I(N__23727));
    LocalMux I__3157 (
            .O(N__23733),
            .I(N__23724));
    Odrv4 I__3156 (
            .O(N__23730),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__3155 (
            .O(N__23727),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv12 I__3154 (
            .O(N__23724),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    CascadeMux I__3153 (
            .O(N__23717),
            .I(N__23714));
    InMux I__3152 (
            .O(N__23714),
            .I(N__23711));
    LocalMux I__3151 (
            .O(N__23711),
            .I(N__23708));
    Odrv4 I__3150 (
            .O(N__23708),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    InMux I__3149 (
            .O(N__23705),
            .I(N__23699));
    InMux I__3148 (
            .O(N__23704),
            .I(N__23695));
    CascadeMux I__3147 (
            .O(N__23703),
            .I(N__23692));
    InMux I__3146 (
            .O(N__23702),
            .I(N__23689));
    LocalMux I__3145 (
            .O(N__23699),
            .I(N__23686));
    InMux I__3144 (
            .O(N__23698),
            .I(N__23683));
    LocalMux I__3143 (
            .O(N__23695),
            .I(N__23680));
    InMux I__3142 (
            .O(N__23692),
            .I(N__23677));
    LocalMux I__3141 (
            .O(N__23689),
            .I(N__23674));
    Span4Mux_h I__3140 (
            .O(N__23686),
            .I(N__23667));
    LocalMux I__3139 (
            .O(N__23683),
            .I(N__23667));
    Span4Mux_v I__3138 (
            .O(N__23680),
            .I(N__23667));
    LocalMux I__3137 (
            .O(N__23677),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv12 I__3136 (
            .O(N__23674),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3135 (
            .O(N__23667),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__3134 (
            .O(N__23660),
            .I(N__23657));
    LocalMux I__3133 (
            .O(N__23657),
            .I(N__23652));
    InMux I__3132 (
            .O(N__23656),
            .I(N__23649));
    CascadeMux I__3131 (
            .O(N__23655),
            .I(N__23645));
    Span4Mux_v I__3130 (
            .O(N__23652),
            .I(N__23641));
    LocalMux I__3129 (
            .O(N__23649),
            .I(N__23638));
    InMux I__3128 (
            .O(N__23648),
            .I(N__23635));
    InMux I__3127 (
            .O(N__23645),
            .I(N__23630));
    InMux I__3126 (
            .O(N__23644),
            .I(N__23630));
    Odrv4 I__3125 (
            .O(N__23641),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3124 (
            .O(N__23638),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3123 (
            .O(N__23635),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3122 (
            .O(N__23630),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__3121 (
            .O(N__23621),
            .I(N__23618));
    InMux I__3120 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__3119 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_h I__3118 (
            .O(N__23612),
            .I(N__23609));
    Odrv4 I__3117 (
            .O(N__23609),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__3116 (
            .O(N__23606),
            .I(N__23603));
    InMux I__3115 (
            .O(N__23603),
            .I(N__23600));
    LocalMux I__3114 (
            .O(N__23600),
            .I(N__23597));
    Span4Mux_h I__3113 (
            .O(N__23597),
            .I(N__23594));
    Odrv4 I__3112 (
            .O(N__23594),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__3111 (
            .O(N__23591),
            .I(N__23587));
    InMux I__3110 (
            .O(N__23590),
            .I(N__23584));
    LocalMux I__3109 (
            .O(N__23587),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__3108 (
            .O(N__23584),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__3107 (
            .O(N__23579),
            .I(N__23576));
    LocalMux I__3106 (
            .O(N__23576),
            .I(N__23571));
    CascadeMux I__3105 (
            .O(N__23575),
            .I(N__23568));
    CascadeMux I__3104 (
            .O(N__23574),
            .I(N__23565));
    Span12Mux_v I__3103 (
            .O(N__23571),
            .I(N__23561));
    InMux I__3102 (
            .O(N__23568),
            .I(N__23558));
    InMux I__3101 (
            .O(N__23565),
            .I(N__23555));
    InMux I__3100 (
            .O(N__23564),
            .I(N__23552));
    Odrv12 I__3099 (
            .O(N__23561),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3098 (
            .O(N__23558),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3097 (
            .O(N__23555),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3096 (
            .O(N__23552),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__3095 (
            .O(N__23543),
            .I(N__23538));
    InMux I__3094 (
            .O(N__23542),
            .I(N__23535));
    InMux I__3093 (
            .O(N__23541),
            .I(N__23532));
    LocalMux I__3092 (
            .O(N__23538),
            .I(N__23527));
    LocalMux I__3091 (
            .O(N__23535),
            .I(N__23527));
    LocalMux I__3090 (
            .O(N__23532),
            .I(N__23524));
    Span4Mux_h I__3089 (
            .O(N__23527),
            .I(N__23521));
    Odrv4 I__3088 (
            .O(N__23524),
            .I(il_min_comp2_D2));
    Odrv4 I__3087 (
            .O(N__23521),
            .I(il_min_comp2_D2));
    InMux I__3086 (
            .O(N__23516),
            .I(N__23511));
    CascadeMux I__3085 (
            .O(N__23515),
            .I(N__23508));
    InMux I__3084 (
            .O(N__23514),
            .I(N__23504));
    LocalMux I__3083 (
            .O(N__23511),
            .I(N__23501));
    InMux I__3082 (
            .O(N__23508),
            .I(N__23496));
    InMux I__3081 (
            .O(N__23507),
            .I(N__23496));
    LocalMux I__3080 (
            .O(N__23504),
            .I(N__23493));
    Span12Mux_v I__3079 (
            .O(N__23501),
            .I(N__23488));
    LocalMux I__3078 (
            .O(N__23496),
            .I(N__23488));
    Odrv4 I__3077 (
            .O(N__23493),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__3076 (
            .O(N__23488),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__3075 (
            .O(N__23483),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__3074 (
            .O(N__23480),
            .I(N__23477));
    LocalMux I__3073 (
            .O(N__23477),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    InMux I__3072 (
            .O(N__23474),
            .I(N__23471));
    LocalMux I__3071 (
            .O(N__23471),
            .I(N__23468));
    Span4Mux_v I__3070 (
            .O(N__23468),
            .I(N__23465));
    Odrv4 I__3069 (
            .O(N__23465),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__3068 (
            .O(N__23462),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ));
    InMux I__3067 (
            .O(N__23459),
            .I(N__23456));
    LocalMux I__3066 (
            .O(N__23456),
            .I(N__23453));
    Odrv4 I__3065 (
            .O(N__23453),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ));
    InMux I__3064 (
            .O(N__23450),
            .I(N__23447));
    LocalMux I__3063 (
            .O(N__23447),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ));
    CascadeMux I__3062 (
            .O(N__23444),
            .I(\delay_measurement_inst.N_30_cascade_ ));
    InMux I__3061 (
            .O(N__23441),
            .I(N__23438));
    LocalMux I__3060 (
            .O(N__23438),
            .I(\delay_measurement_inst.N_37 ));
    IoInMux I__3059 (
            .O(N__23435),
            .I(N__23432));
    LocalMux I__3058 (
            .O(N__23432),
            .I(N__23429));
    Span4Mux_s3_v I__3057 (
            .O(N__23429),
            .I(N__23426));
    Span4Mux_v I__3056 (
            .O(N__23426),
            .I(N__23423));
    Odrv4 I__3055 (
            .O(N__23423),
            .I(\delay_measurement_inst.delay_hc_timer.N_302_i ));
    InMux I__3054 (
            .O(N__23420),
            .I(N__23417));
    LocalMux I__3053 (
            .O(N__23417),
            .I(\delay_measurement_inst.N_36 ));
    InMux I__3052 (
            .O(N__23414),
            .I(N__23411));
    LocalMux I__3051 (
            .O(N__23411),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    CascadeMux I__3050 (
            .O(N__23408),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9_cascade_ ));
    CascadeMux I__3049 (
            .O(N__23405),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_ ));
    InMux I__3048 (
            .O(N__23402),
            .I(N__23399));
    LocalMux I__3047 (
            .O(N__23399),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ));
    CascadeMux I__3046 (
            .O(N__23396),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12_cascade_ ));
    InMux I__3045 (
            .O(N__23393),
            .I(N__23390));
    LocalMux I__3044 (
            .O(N__23390),
            .I(N__23387));
    Odrv12 I__3043 (
            .O(N__23387),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ));
    CascadeMux I__3042 (
            .O(N__23384),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_4_cascade_ ));
    InMux I__3041 (
            .O(N__23381),
            .I(N__23378));
    LocalMux I__3040 (
            .O(N__23378),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0 ));
    CascadeMux I__3039 (
            .O(N__23375),
            .I(\delay_measurement_inst.un1_elapsed_time_hc_cascade_ ));
    InMux I__3038 (
            .O(N__23372),
            .I(N__23369));
    LocalMux I__3037 (
            .O(N__23369),
            .I(\delay_measurement_inst.N_31 ));
    InMux I__3036 (
            .O(N__23366),
            .I(N__23363));
    LocalMux I__3035 (
            .O(N__23363),
            .I(\delay_measurement_inst.N_40 ));
    InMux I__3034 (
            .O(N__23360),
            .I(N__23357));
    LocalMux I__3033 (
            .O(N__23357),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ));
    CascadeMux I__3032 (
            .O(N__23354),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_ ));
    InMux I__3031 (
            .O(N__23351),
            .I(N__23348));
    LocalMux I__3030 (
            .O(N__23348),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8 ));
    CascadeMux I__3029 (
            .O(N__23345),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1_cascade_ ));
    InMux I__3028 (
            .O(N__23342),
            .I(N__23339));
    LocalMux I__3027 (
            .O(N__23339),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt14_0 ));
    CascadeMux I__3026 (
            .O(N__23336),
            .I(N__23333));
    InMux I__3025 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__3024 (
            .O(N__23330),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__3023 (
            .O(N__23327),
            .I(N__23324));
    InMux I__3022 (
            .O(N__23324),
            .I(N__23321));
    LocalMux I__3021 (
            .O(N__23321),
            .I(N__23318));
    Odrv4 I__3020 (
            .O(N__23318),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__3019 (
            .O(N__23315),
            .I(N__23312));
    InMux I__3018 (
            .O(N__23312),
            .I(N__23309));
    LocalMux I__3017 (
            .O(N__23309),
            .I(N__23306));
    Odrv4 I__3016 (
            .O(N__23306),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__3015 (
            .O(N__23303),
            .I(N__23300));
    InMux I__3014 (
            .O(N__23300),
            .I(N__23297));
    LocalMux I__3013 (
            .O(N__23297),
            .I(N__23294));
    Span4Mux_h I__3012 (
            .O(N__23294),
            .I(N__23291));
    Odrv4 I__3011 (
            .O(N__23291),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__3010 (
            .O(N__23288),
            .I(N__23285));
    InMux I__3009 (
            .O(N__23285),
            .I(N__23282));
    LocalMux I__3008 (
            .O(N__23282),
            .I(N__23279));
    Span4Mux_v I__3007 (
            .O(N__23279),
            .I(N__23276));
    Odrv4 I__3006 (
            .O(N__23276),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__3005 (
            .O(N__23273),
            .I(N__23270));
    InMux I__3004 (
            .O(N__23270),
            .I(N__23267));
    LocalMux I__3003 (
            .O(N__23267),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__3002 (
            .O(N__23264),
            .I(N__23261));
    InMux I__3001 (
            .O(N__23261),
            .I(N__23258));
    LocalMux I__3000 (
            .O(N__23258),
            .I(N__23255));
    Span4Mux_v I__2999 (
            .O(N__23255),
            .I(N__23252));
    Odrv4 I__2998 (
            .O(N__23252),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    IoInMux I__2997 (
            .O(N__23249),
            .I(N__23246));
    LocalMux I__2996 (
            .O(N__23246),
            .I(N__23243));
    Span12Mux_s8_v I__2995 (
            .O(N__23243),
            .I(N__23240));
    Odrv12 I__2994 (
            .O(N__23240),
            .I(s4_phy_c));
    CascadeMux I__2993 (
            .O(N__23237),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__2992 (
            .O(N__23234),
            .I(N__23231));
    InMux I__2991 (
            .O(N__23231),
            .I(N__23228));
    LocalMux I__2990 (
            .O(N__23228),
            .I(N__23225));
    Odrv4 I__2989 (
            .O(N__23225),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__2988 (
            .O(N__23222),
            .I(N__23219));
    InMux I__2987 (
            .O(N__23219),
            .I(N__23216));
    LocalMux I__2986 (
            .O(N__23216),
            .I(N__23213));
    Odrv12 I__2985 (
            .O(N__23213),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    InMux I__2984 (
            .O(N__23210),
            .I(N__23207));
    LocalMux I__2983 (
            .O(N__23207),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__2982 (
            .O(N__23204),
            .I(N__23201));
    LocalMux I__2981 (
            .O(N__23201),
            .I(N__23198));
    Span4Mux_v I__2980 (
            .O(N__23198),
            .I(N__23195));
    Odrv4 I__2979 (
            .O(N__23195),
            .I(\current_shift_inst.PI_CTRL.N_71 ));
    CascadeMux I__2978 (
            .O(N__23192),
            .I(\current_shift_inst.PI_CTRL.N_75_cascade_ ));
    CascadeMux I__2977 (
            .O(N__23189),
            .I(N__23186));
    InMux I__2976 (
            .O(N__23186),
            .I(N__23183));
    LocalMux I__2975 (
            .O(N__23183),
            .I(N__23180));
    Odrv4 I__2974 (
            .O(N__23180),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    CascadeMux I__2973 (
            .O(N__23177),
            .I(N__23174));
    InMux I__2972 (
            .O(N__23174),
            .I(N__23171));
    LocalMux I__2971 (
            .O(N__23171),
            .I(N__23168));
    Span4Mux_v I__2970 (
            .O(N__23168),
            .I(N__23165));
    Odrv4 I__2969 (
            .O(N__23165),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__2968 (
            .O(N__23162),
            .I(N__23159));
    InMux I__2967 (
            .O(N__23159),
            .I(N__23156));
    LocalMux I__2966 (
            .O(N__23156),
            .I(N__23153));
    Odrv4 I__2965 (
            .O(N__23153),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__2964 (
            .O(N__23150),
            .I(N__23147));
    InMux I__2963 (
            .O(N__23147),
            .I(N__23144));
    LocalMux I__2962 (
            .O(N__23144),
            .I(N__23141));
    Odrv4 I__2961 (
            .O(N__23141),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__2960 (
            .O(N__23138),
            .I(N__23135));
    LocalMux I__2959 (
            .O(N__23135),
            .I(N__23132));
    Odrv4 I__2958 (
            .O(N__23132),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    InMux I__2957 (
            .O(N__23129),
            .I(N__23126));
    LocalMux I__2956 (
            .O(N__23126),
            .I(N__23123));
    Odrv4 I__2955 (
            .O(N__23123),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__2954 (
            .O(N__23120),
            .I(N__23117));
    LocalMux I__2953 (
            .O(N__23117),
            .I(N__23114));
    Odrv4 I__2952 (
            .O(N__23114),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    CascadeMux I__2951 (
            .O(N__23111),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ));
    CascadeMux I__2950 (
            .O(N__23108),
            .I(\current_shift_inst.PI_CTRL.N_74_cascade_ ));
    InMux I__2949 (
            .O(N__23105),
            .I(N__23102));
    LocalMux I__2948 (
            .O(N__23102),
            .I(N__23099));
    Odrv4 I__2947 (
            .O(N__23099),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__2946 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__2945 (
            .O(N__23093),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    CascadeMux I__2944 (
            .O(N__23090),
            .I(N__23087));
    InMux I__2943 (
            .O(N__23087),
            .I(N__23084));
    LocalMux I__2942 (
            .O(N__23084),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    InMux I__2941 (
            .O(N__23081),
            .I(N__23078));
    LocalMux I__2940 (
            .O(N__23078),
            .I(\delay_measurement_inst.N_32 ));
    InMux I__2939 (
            .O(N__23075),
            .I(N__23072));
    LocalMux I__2938 (
            .O(N__23072),
            .I(\delay_measurement_inst.N_35 ));
    InMux I__2937 (
            .O(N__23069),
            .I(N__23066));
    LocalMux I__2936 (
            .O(N__23066),
            .I(N__23063));
    Odrv4 I__2935 (
            .O(N__23063),
            .I(\delay_measurement_inst.N_43 ));
    InMux I__2934 (
            .O(N__23060),
            .I(N__23057));
    LocalMux I__2933 (
            .O(N__23057),
            .I(N__23054));
    Odrv12 I__2932 (
            .O(N__23054),
            .I(il_max_comp1_c));
    InMux I__2931 (
            .O(N__23051),
            .I(N__23048));
    LocalMux I__2930 (
            .O(N__23048),
            .I(N__23045));
    Span4Mux_v I__2929 (
            .O(N__23045),
            .I(N__23042));
    Odrv4 I__2928 (
            .O(N__23042),
            .I(\delay_measurement_inst.N_34 ));
    CascadeMux I__2927 (
            .O(N__23039),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_ ));
    InMux I__2926 (
            .O(N__23036),
            .I(N__23033));
    LocalMux I__2925 (
            .O(N__23033),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__2924 (
            .O(N__23030),
            .I(N__23027));
    LocalMux I__2923 (
            .O(N__23027),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__2922 (
            .O(N__23024),
            .I(N__23021));
    LocalMux I__2921 (
            .O(N__23021),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__2920 (
            .O(N__23018),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__2919 (
            .O(N__23015),
            .I(N__23012));
    InMux I__2918 (
            .O(N__23012),
            .I(N__23009));
    LocalMux I__2917 (
            .O(N__23009),
            .I(N__23006));
    Odrv4 I__2916 (
            .O(N__23006),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__2915 (
            .O(N__23003),
            .I(N__23000));
    InMux I__2914 (
            .O(N__23000),
            .I(N__22997));
    LocalMux I__2913 (
            .O(N__22997),
            .I(N__22994));
    Odrv4 I__2912 (
            .O(N__22994),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__2911 (
            .O(N__22991),
            .I(N__22988));
    InMux I__2910 (
            .O(N__22988),
            .I(N__22985));
    LocalMux I__2909 (
            .O(N__22985),
            .I(N__22982));
    Span4Mux_h I__2908 (
            .O(N__22982),
            .I(N__22979));
    Odrv4 I__2907 (
            .O(N__22979),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__2906 (
            .O(N__22976),
            .I(N__22973));
    InMux I__2905 (
            .O(N__22973),
            .I(N__22970));
    LocalMux I__2904 (
            .O(N__22970),
            .I(N__22967));
    Odrv12 I__2903 (
            .O(N__22967),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    InMux I__2902 (
            .O(N__22964),
            .I(N__22961));
    LocalMux I__2901 (
            .O(N__22961),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__2900 (
            .O(N__22958),
            .I(N__22955));
    InMux I__2899 (
            .O(N__22955),
            .I(N__22952));
    LocalMux I__2898 (
            .O(N__22952),
            .I(N__22949));
    Span4Mux_h I__2897 (
            .O(N__22949),
            .I(N__22946));
    Span4Mux_h I__2896 (
            .O(N__22946),
            .I(N__22943));
    Odrv4 I__2895 (
            .O(N__22943),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__2894 (
            .O(N__22940),
            .I(N__22937));
    LocalMux I__2893 (
            .O(N__22937),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__2892 (
            .O(N__22934),
            .I(N__22931));
    InMux I__2891 (
            .O(N__22931),
            .I(N__22928));
    LocalMux I__2890 (
            .O(N__22928),
            .I(N__22925));
    Span4Mux_h I__2889 (
            .O(N__22925),
            .I(N__22922));
    Span4Mux_h I__2888 (
            .O(N__22922),
            .I(N__22919));
    Odrv4 I__2887 (
            .O(N__22919),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__2886 (
            .O(N__22916),
            .I(N__22913));
    LocalMux I__2885 (
            .O(N__22913),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__2884 (
            .O(N__22910),
            .I(N__22907));
    LocalMux I__2883 (
            .O(N__22907),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__2882 (
            .O(N__22904),
            .I(N__22901));
    LocalMux I__2881 (
            .O(N__22901),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__2880 (
            .O(N__22898),
            .I(N__22895));
    LocalMux I__2879 (
            .O(N__22895),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__2878 (
            .O(N__22892),
            .I(N__22889));
    LocalMux I__2877 (
            .O(N__22889),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__2876 (
            .O(N__22886),
            .I(N__22883));
    LocalMux I__2875 (
            .O(N__22883),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__2874 (
            .O(N__22880),
            .I(N__22877));
    LocalMux I__2873 (
            .O(N__22877),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__2872 (
            .O(N__22874),
            .I(N__22871));
    LocalMux I__2871 (
            .O(N__22871),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__2870 (
            .O(N__22868),
            .I(N__22865));
    LocalMux I__2869 (
            .O(N__22865),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__2868 (
            .O(N__22862),
            .I(N__22859));
    LocalMux I__2867 (
            .O(N__22859),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__2866 (
            .O(N__22856),
            .I(N__22853));
    LocalMux I__2865 (
            .O(N__22853),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__2864 (
            .O(N__22850),
            .I(N__22847));
    LocalMux I__2863 (
            .O(N__22847),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__2862 (
            .O(N__22844),
            .I(N__22841));
    LocalMux I__2861 (
            .O(N__22841),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__2860 (
            .O(N__22838),
            .I(N__22835));
    LocalMux I__2859 (
            .O(N__22835),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__2858 (
            .O(N__22832),
            .I(N__22826));
    InMux I__2857 (
            .O(N__22831),
            .I(N__22826));
    LocalMux I__2856 (
            .O(N__22826),
            .I(N__22823));
    Odrv4 I__2855 (
            .O(N__22823),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2854 (
            .O(N__22820),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__2853 (
            .O(N__22817),
            .I(N__22811));
    InMux I__2852 (
            .O(N__22816),
            .I(N__22811));
    LocalMux I__2851 (
            .O(N__22811),
            .I(N__22808));
    Odrv4 I__2850 (
            .O(N__22808),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2849 (
            .O(N__22805),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2848 (
            .O(N__22802),
            .I(N__22796));
    InMux I__2847 (
            .O(N__22801),
            .I(N__22796));
    LocalMux I__2846 (
            .O(N__22796),
            .I(N__22793));
    Odrv4 I__2845 (
            .O(N__22793),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2844 (
            .O(N__22790),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2843 (
            .O(N__22787),
            .I(N__22783));
    InMux I__2842 (
            .O(N__22786),
            .I(N__22780));
    LocalMux I__2841 (
            .O(N__22783),
            .I(N__22775));
    LocalMux I__2840 (
            .O(N__22780),
            .I(N__22775));
    Span4Mux_h I__2839 (
            .O(N__22775),
            .I(N__22772));
    Odrv4 I__2838 (
            .O(N__22772),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2837 (
            .O(N__22769),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2836 (
            .O(N__22766),
            .I(N__22763));
    LocalMux I__2835 (
            .O(N__22763),
            .I(N__22759));
    InMux I__2834 (
            .O(N__22762),
            .I(N__22756));
    Span4Mux_h I__2833 (
            .O(N__22759),
            .I(N__22751));
    LocalMux I__2832 (
            .O(N__22756),
            .I(N__22751));
    Odrv4 I__2831 (
            .O(N__22751),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2830 (
            .O(N__22748),
            .I(bfn_7_14_0_));
    InMux I__2829 (
            .O(N__22745),
            .I(N__22742));
    LocalMux I__2828 (
            .O(N__22742),
            .I(N__22738));
    InMux I__2827 (
            .O(N__22741),
            .I(N__22735));
    Span4Mux_v I__2826 (
            .O(N__22738),
            .I(N__22732));
    LocalMux I__2825 (
            .O(N__22735),
            .I(N__22729));
    Odrv4 I__2824 (
            .O(N__22732),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    Odrv12 I__2823 (
            .O(N__22729),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2822 (
            .O(N__22724),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2821 (
            .O(N__22721),
            .I(N__22717));
    InMux I__2820 (
            .O(N__22720),
            .I(N__22714));
    LocalMux I__2819 (
            .O(N__22717),
            .I(N__22709));
    LocalMux I__2818 (
            .O(N__22714),
            .I(N__22709));
    Odrv4 I__2817 (
            .O(N__22709),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2816 (
            .O(N__22706),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2815 (
            .O(N__22703),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2814 (
            .O(N__22700),
            .I(N__22696));
    CascadeMux I__2813 (
            .O(N__22699),
            .I(N__22693));
    LocalMux I__2812 (
            .O(N__22696),
            .I(N__22686));
    InMux I__2811 (
            .O(N__22693),
            .I(N__22683));
    CascadeMux I__2810 (
            .O(N__22692),
            .I(N__22680));
    CascadeMux I__2809 (
            .O(N__22691),
            .I(N__22677));
    CascadeMux I__2808 (
            .O(N__22690),
            .I(N__22674));
    CascadeMux I__2807 (
            .O(N__22689),
            .I(N__22670));
    Span4Mux_s2_h I__2806 (
            .O(N__22686),
            .I(N__22662));
    LocalMux I__2805 (
            .O(N__22683),
            .I(N__22662));
    InMux I__2804 (
            .O(N__22680),
            .I(N__22655));
    InMux I__2803 (
            .O(N__22677),
            .I(N__22655));
    InMux I__2802 (
            .O(N__22674),
            .I(N__22655));
    InMux I__2801 (
            .O(N__22673),
            .I(N__22652));
    InMux I__2800 (
            .O(N__22670),
            .I(N__22649));
    InMux I__2799 (
            .O(N__22669),
            .I(N__22646));
    InMux I__2798 (
            .O(N__22668),
            .I(N__22641));
    InMux I__2797 (
            .O(N__22667),
            .I(N__22641));
    Span4Mux_v I__2796 (
            .O(N__22662),
            .I(N__22638));
    LocalMux I__2795 (
            .O(N__22655),
            .I(N__22633));
    LocalMux I__2794 (
            .O(N__22652),
            .I(N__22633));
    LocalMux I__2793 (
            .O(N__22649),
            .I(N__22626));
    LocalMux I__2792 (
            .O(N__22646),
            .I(N__22626));
    LocalMux I__2791 (
            .O(N__22641),
            .I(N__22626));
    Span4Mux_v I__2790 (
            .O(N__22638),
            .I(N__22623));
    Span4Mux_s3_h I__2789 (
            .O(N__22633),
            .I(N__22620));
    Span4Mux_h I__2788 (
            .O(N__22626),
            .I(N__22617));
    Span4Mux_h I__2787 (
            .O(N__22623),
            .I(N__22614));
    Span4Mux_h I__2786 (
            .O(N__22620),
            .I(N__22611));
    Span4Mux_h I__2785 (
            .O(N__22617),
            .I(N__22608));
    Odrv4 I__2784 (
            .O(N__22614),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2783 (
            .O(N__22611),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2782 (
            .O(N__22608),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__2781 (
            .O(N__22601),
            .I(N__22598));
    InMux I__2780 (
            .O(N__22598),
            .I(N__22594));
    CascadeMux I__2779 (
            .O(N__22597),
            .I(N__22591));
    LocalMux I__2778 (
            .O(N__22594),
            .I(N__22588));
    InMux I__2777 (
            .O(N__22591),
            .I(N__22585));
    Span4Mux_v I__2776 (
            .O(N__22588),
            .I(N__22580));
    LocalMux I__2775 (
            .O(N__22585),
            .I(N__22580));
    Odrv4 I__2774 (
            .O(N__22580),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2773 (
            .O(N__22577),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__2772 (
            .O(N__22574),
            .I(N__22568));
    InMux I__2771 (
            .O(N__22573),
            .I(N__22568));
    LocalMux I__2770 (
            .O(N__22568),
            .I(N__22565));
    Odrv4 I__2769 (
            .O(N__22565),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2768 (
            .O(N__22562),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2767 (
            .O(N__22559),
            .I(N__22553));
    InMux I__2766 (
            .O(N__22558),
            .I(N__22553));
    LocalMux I__2765 (
            .O(N__22553),
            .I(N__22550));
    Span4Mux_v I__2764 (
            .O(N__22550),
            .I(N__22547));
    Odrv4 I__2763 (
            .O(N__22547),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2762 (
            .O(N__22544),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2761 (
            .O(N__22541),
            .I(N__22538));
    LocalMux I__2760 (
            .O(N__22538),
            .I(N__22534));
    InMux I__2759 (
            .O(N__22537),
            .I(N__22531));
    Span4Mux_v I__2758 (
            .O(N__22534),
            .I(N__22526));
    LocalMux I__2757 (
            .O(N__22531),
            .I(N__22526));
    Odrv4 I__2756 (
            .O(N__22526),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2755 (
            .O(N__22523),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2754 (
            .O(N__22520),
            .I(N__22516));
    InMux I__2753 (
            .O(N__22519),
            .I(N__22513));
    LocalMux I__2752 (
            .O(N__22516),
            .I(N__22510));
    LocalMux I__2751 (
            .O(N__22513),
            .I(N__22507));
    Span4Mux_h I__2750 (
            .O(N__22510),
            .I(N__22502));
    Span4Mux_v I__2749 (
            .O(N__22507),
            .I(N__22502));
    Odrv4 I__2748 (
            .O(N__22502),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2747 (
            .O(N__22499),
            .I(bfn_7_13_0_));
    InMux I__2746 (
            .O(N__22496),
            .I(N__22490));
    InMux I__2745 (
            .O(N__22495),
            .I(N__22490));
    LocalMux I__2744 (
            .O(N__22490),
            .I(N__22487));
    Odrv4 I__2743 (
            .O(N__22487),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2742 (
            .O(N__22484),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__2741 (
            .O(N__22481),
            .I(N__22478));
    InMux I__2740 (
            .O(N__22478),
            .I(N__22472));
    InMux I__2739 (
            .O(N__22477),
            .I(N__22472));
    LocalMux I__2738 (
            .O(N__22472),
            .I(N__22469));
    Span4Mux_h I__2737 (
            .O(N__22469),
            .I(N__22466));
    Odrv4 I__2736 (
            .O(N__22466),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2735 (
            .O(N__22463),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__2734 (
            .O(N__22460),
            .I(N__22456));
    InMux I__2733 (
            .O(N__22459),
            .I(N__22453));
    InMux I__2732 (
            .O(N__22456),
            .I(N__22450));
    LocalMux I__2731 (
            .O(N__22453),
            .I(N__22445));
    LocalMux I__2730 (
            .O(N__22450),
            .I(N__22445));
    Odrv4 I__2729 (
            .O(N__22445),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2728 (
            .O(N__22442),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2727 (
            .O(N__22439),
            .I(N__22436));
    InMux I__2726 (
            .O(N__22436),
            .I(N__22433));
    LocalMux I__2725 (
            .O(N__22433),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__2724 (
            .O(N__22430),
            .I(N__22425));
    InMux I__2723 (
            .O(N__22429),
            .I(N__22420));
    InMux I__2722 (
            .O(N__22428),
            .I(N__22420));
    LocalMux I__2721 (
            .O(N__22425),
            .I(N__22415));
    LocalMux I__2720 (
            .O(N__22420),
            .I(N__22415));
    Odrv12 I__2719 (
            .O(N__22415),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2718 (
            .O(N__22412),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    CascadeMux I__2717 (
            .O(N__22409),
            .I(N__22406));
    InMux I__2716 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__2715 (
            .O(N__22403),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2714 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__2713 (
            .O(N__22397),
            .I(N__22394));
    Span4Mux_v I__2712 (
            .O(N__22394),
            .I(N__22389));
    InMux I__2711 (
            .O(N__22393),
            .I(N__22384));
    InMux I__2710 (
            .O(N__22392),
            .I(N__22384));
    Sp12to4 I__2709 (
            .O(N__22389),
            .I(N__22379));
    LocalMux I__2708 (
            .O(N__22384),
            .I(N__22379));
    Odrv12 I__2707 (
            .O(N__22379),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2706 (
            .O(N__22376),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    CascadeMux I__2705 (
            .O(N__22373),
            .I(N__22370));
    InMux I__2704 (
            .O(N__22370),
            .I(N__22367));
    LocalMux I__2703 (
            .O(N__22367),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2702 (
            .O(N__22364),
            .I(N__22360));
    InMux I__2701 (
            .O(N__22363),
            .I(N__22357));
    LocalMux I__2700 (
            .O(N__22360),
            .I(N__22354));
    LocalMux I__2699 (
            .O(N__22357),
            .I(N__22351));
    Span4Mux_h I__2698 (
            .O(N__22354),
            .I(N__22348));
    Span4Mux_h I__2697 (
            .O(N__22351),
            .I(N__22345));
    Odrv4 I__2696 (
            .O(N__22348),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    Odrv4 I__2695 (
            .O(N__22345),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2694 (
            .O(N__22340),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    CascadeMux I__2693 (
            .O(N__22337),
            .I(N__22333));
    CascadeMux I__2692 (
            .O(N__22336),
            .I(N__22330));
    InMux I__2691 (
            .O(N__22333),
            .I(N__22327));
    InMux I__2690 (
            .O(N__22330),
            .I(N__22324));
    LocalMux I__2689 (
            .O(N__22327),
            .I(N__22321));
    LocalMux I__2688 (
            .O(N__22324),
            .I(N__22318));
    Span4Mux_h I__2687 (
            .O(N__22321),
            .I(N__22315));
    Span4Mux_h I__2686 (
            .O(N__22318),
            .I(N__22312));
    Odrv4 I__2685 (
            .O(N__22315),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    Odrv4 I__2684 (
            .O(N__22312),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2683 (
            .O(N__22307),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2682 (
            .O(N__22304),
            .I(N__22301));
    LocalMux I__2681 (
            .O(N__22301),
            .I(N__22298));
    Odrv4 I__2680 (
            .O(N__22298),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2679 (
            .O(N__22295),
            .I(N__22291));
    InMux I__2678 (
            .O(N__22294),
            .I(N__22288));
    LocalMux I__2677 (
            .O(N__22291),
            .I(N__22285));
    LocalMux I__2676 (
            .O(N__22288),
            .I(N__22282));
    Span4Mux_h I__2675 (
            .O(N__22285),
            .I(N__22279));
    Odrv12 I__2674 (
            .O(N__22282),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    Odrv4 I__2673 (
            .O(N__22279),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2672 (
            .O(N__22274),
            .I(bfn_7_12_0_));
    InMux I__2671 (
            .O(N__22271),
            .I(N__22265));
    InMux I__2670 (
            .O(N__22270),
            .I(N__22265));
    LocalMux I__2669 (
            .O(N__22265),
            .I(N__22262));
    Odrv4 I__2668 (
            .O(N__22262),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2667 (
            .O(N__22259),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2666 (
            .O(N__22256),
            .I(N__22250));
    InMux I__2665 (
            .O(N__22255),
            .I(N__22250));
    LocalMux I__2664 (
            .O(N__22250),
            .I(N__22247));
    Odrv4 I__2663 (
            .O(N__22247),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2662 (
            .O(N__22244),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2661 (
            .O(N__22241),
            .I(N__22235));
    InMux I__2660 (
            .O(N__22240),
            .I(N__22235));
    LocalMux I__2659 (
            .O(N__22235),
            .I(N__22232));
    Odrv4 I__2658 (
            .O(N__22232),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2657 (
            .O(N__22229),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2656 (
            .O(N__22226),
            .I(N__22223));
    InMux I__2655 (
            .O(N__22223),
            .I(N__22220));
    LocalMux I__2654 (
            .O(N__22220),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2653 (
            .O(N__22217),
            .I(N__22213));
    CascadeMux I__2652 (
            .O(N__22216),
            .I(N__22210));
    InMux I__2651 (
            .O(N__22213),
            .I(N__22205));
    InMux I__2650 (
            .O(N__22210),
            .I(N__22198));
    InMux I__2649 (
            .O(N__22209),
            .I(N__22198));
    InMux I__2648 (
            .O(N__22208),
            .I(N__22198));
    LocalMux I__2647 (
            .O(N__22205),
            .I(N__22195));
    LocalMux I__2646 (
            .O(N__22198),
            .I(N__22192));
    Span4Mux_v I__2645 (
            .O(N__22195),
            .I(N__22187));
    Span4Mux_v I__2644 (
            .O(N__22192),
            .I(N__22187));
    Span4Mux_h I__2643 (
            .O(N__22187),
            .I(N__22184));
    Odrv4 I__2642 (
            .O(N__22184),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2641 (
            .O(N__22181),
            .I(N__22178));
    LocalMux I__2640 (
            .O(N__22178),
            .I(N__22173));
    InMux I__2639 (
            .O(N__22177),
            .I(N__22168));
    InMux I__2638 (
            .O(N__22176),
            .I(N__22168));
    Span12Mux_s2_h I__2637 (
            .O(N__22173),
            .I(N__22163));
    LocalMux I__2636 (
            .O(N__22168),
            .I(N__22163));
    Odrv12 I__2635 (
            .O(N__22163),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2634 (
            .O(N__22160),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2633 (
            .O(N__22157),
            .I(N__22152));
    InMux I__2632 (
            .O(N__22156),
            .I(N__22147));
    InMux I__2631 (
            .O(N__22155),
            .I(N__22147));
    LocalMux I__2630 (
            .O(N__22152),
            .I(N__22142));
    LocalMux I__2629 (
            .O(N__22147),
            .I(N__22142));
    Odrv12 I__2628 (
            .O(N__22142),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2627 (
            .O(N__22139),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2626 (
            .O(N__22136),
            .I(N__22133));
    LocalMux I__2625 (
            .O(N__22133),
            .I(N__22128));
    InMux I__2624 (
            .O(N__22132),
            .I(N__22123));
    InMux I__2623 (
            .O(N__22131),
            .I(N__22123));
    Span12Mux_s7_h I__2622 (
            .O(N__22128),
            .I(N__22120));
    LocalMux I__2621 (
            .O(N__22123),
            .I(N__22117));
    Odrv12 I__2620 (
            .O(N__22120),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv12 I__2619 (
            .O(N__22117),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2618 (
            .O(N__22112),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2617 (
            .O(N__22109),
            .I(N__22106));
    LocalMux I__2616 (
            .O(N__22106),
            .I(N__22103));
    Odrv4 I__2615 (
            .O(N__22103),
            .I(il_min_comp2_c));
    InMux I__2614 (
            .O(N__22100),
            .I(N__22097));
    LocalMux I__2613 (
            .O(N__22097),
            .I(N__22094));
    Odrv4 I__2612 (
            .O(N__22094),
            .I(il_min_comp2_D1));
    CascadeMux I__2611 (
            .O(N__22091),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    CascadeMux I__2610 (
            .O(N__22088),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ));
    CascadeMux I__2609 (
            .O(N__22085),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    CascadeMux I__2608 (
            .O(N__22082),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2607 (
            .O(N__22079),
            .I(N__22076));
    LocalMux I__2606 (
            .O(N__22076),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2605 (
            .O(N__22073),
            .I(N__22070));
    LocalMux I__2604 (
            .O(N__22070),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2603 (
            .O(N__22067),
            .I(N__22064));
    LocalMux I__2602 (
            .O(N__22064),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2601 (
            .O(N__22061),
            .I(N__22058));
    LocalMux I__2600 (
            .O(N__22058),
            .I(N__22055));
    Odrv4 I__2599 (
            .O(N__22055),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__2598 (
            .O(N__22052),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ));
    InMux I__2597 (
            .O(N__22049),
            .I(N__22046));
    LocalMux I__2596 (
            .O(N__22046),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2595 (
            .O(N__22043),
            .I(N__22040));
    LocalMux I__2594 (
            .O(N__22040),
            .I(N__22031));
    InMux I__2593 (
            .O(N__22039),
            .I(N__22024));
    InMux I__2592 (
            .O(N__22038),
            .I(N__22024));
    InMux I__2591 (
            .O(N__22037),
            .I(N__22024));
    InMux I__2590 (
            .O(N__22036),
            .I(N__22019));
    InMux I__2589 (
            .O(N__22035),
            .I(N__22019));
    InMux I__2588 (
            .O(N__22034),
            .I(N__22016));
    Span4Mux_v I__2587 (
            .O(N__22031),
            .I(N__22011));
    LocalMux I__2586 (
            .O(N__22024),
            .I(N__22011));
    LocalMux I__2585 (
            .O(N__22019),
            .I(N__22006));
    LocalMux I__2584 (
            .O(N__22016),
            .I(N__22006));
    Span4Mux_h I__2583 (
            .O(N__22011),
            .I(N__22003));
    Span4Mux_h I__2582 (
            .O(N__22006),
            .I(N__22000));
    Odrv4 I__2581 (
            .O(N__22003),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2580 (
            .O(N__22000),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2579 (
            .O(N__21995),
            .I(N__21992));
    LocalMux I__2578 (
            .O(N__21992),
            .I(N__21989));
    Span4Mux_v I__2577 (
            .O(N__21989),
            .I(N__21986));
    Odrv4 I__2576 (
            .O(N__21986),
            .I(il_max_comp2_D1));
    InMux I__2575 (
            .O(N__21983),
            .I(N__21980));
    LocalMux I__2574 (
            .O(N__21980),
            .I(N__21977));
    Odrv12 I__2573 (
            .O(N__21977),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2572 (
            .O(N__21974),
            .I(N__21971));
    LocalMux I__2571 (
            .O(N__21971),
            .I(N__21968));
    Span4Mux_s3_h I__2570 (
            .O(N__21968),
            .I(N__21965));
    Odrv4 I__2569 (
            .O(N__21965),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2568 (
            .O(N__21962),
            .I(N__21959));
    LocalMux I__2567 (
            .O(N__21959),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2566 (
            .O(N__21956),
            .I(N__21953));
    InMux I__2565 (
            .O(N__21953),
            .I(N__21950));
    LocalMux I__2564 (
            .O(N__21950),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2563 (
            .O(N__21947),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__2562 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__2561 (
            .O(N__21941),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    CascadeMux I__2560 (
            .O(N__21938),
            .I(N__21935));
    InMux I__2559 (
            .O(N__21935),
            .I(N__21932));
    LocalMux I__2558 (
            .O(N__21932),
            .I(N__21929));
    Span4Mux_v I__2557 (
            .O(N__21929),
            .I(N__21926));
    Odrv4 I__2556 (
            .O(N__21926),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2555 (
            .O(N__21923),
            .I(N__21918));
    InMux I__2554 (
            .O(N__21922),
            .I(N__21915));
    InMux I__2553 (
            .O(N__21921),
            .I(N__21912));
    LocalMux I__2552 (
            .O(N__21918),
            .I(N__21909));
    LocalMux I__2551 (
            .O(N__21915),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2550 (
            .O(N__21912),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2549 (
            .O(N__21909),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2548 (
            .O(N__21902),
            .I(N__21899));
    LocalMux I__2547 (
            .O(N__21899),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2546 (
            .O(N__21896),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2545 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__2544 (
            .O(N__21890),
            .I(N__21887));
    Span12Mux_s9_v I__2543 (
            .O(N__21887),
            .I(N__21884));
    Span12Mux_h I__2542 (
            .O(N__21884),
            .I(N__21881));
    Odrv12 I__2541 (
            .O(N__21881),
            .I(pwm_output_c));
    CascadeMux I__2540 (
            .O(N__21878),
            .I(N__21874));
    InMux I__2539 (
            .O(N__21877),
            .I(N__21864));
    InMux I__2538 (
            .O(N__21874),
            .I(N__21859));
    InMux I__2537 (
            .O(N__21873),
            .I(N__21859));
    InMux I__2536 (
            .O(N__21872),
            .I(N__21854));
    InMux I__2535 (
            .O(N__21871),
            .I(N__21854));
    InMux I__2534 (
            .O(N__21870),
            .I(N__21847));
    InMux I__2533 (
            .O(N__21869),
            .I(N__21847));
    InMux I__2532 (
            .O(N__21868),
            .I(N__21847));
    InMux I__2531 (
            .O(N__21867),
            .I(N__21844));
    LocalMux I__2530 (
            .O(N__21864),
            .I(N__21841));
    LocalMux I__2529 (
            .O(N__21859),
            .I(N__21836));
    LocalMux I__2528 (
            .O(N__21854),
            .I(N__21836));
    LocalMux I__2527 (
            .O(N__21847),
            .I(N__21831));
    LocalMux I__2526 (
            .O(N__21844),
            .I(N__21831));
    Span4Mux_h I__2525 (
            .O(N__21841),
            .I(N__21828));
    Span4Mux_h I__2524 (
            .O(N__21836),
            .I(N__21825));
    Span4Mux_h I__2523 (
            .O(N__21831),
            .I(N__21822));
    Odrv4 I__2522 (
            .O(N__21828),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2521 (
            .O(N__21825),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2520 (
            .O(N__21822),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    CascadeMux I__2519 (
            .O(N__21815),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__2518 (
            .O(N__21812),
            .I(N__21809));
    LocalMux I__2517 (
            .O(N__21809),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2516 (
            .O(N__21806),
            .I(N__21803));
    LocalMux I__2515 (
            .O(N__21803),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    CascadeMux I__2514 (
            .O(N__21800),
            .I(N__21797));
    InMux I__2513 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__2512 (
            .O(N__21794),
            .I(N__21791));
    Odrv12 I__2511 (
            .O(N__21791),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__2510 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__2509 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__2508 (
            .O(N__21782),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    CascadeMux I__2507 (
            .O(N__21779),
            .I(N__21776));
    InMux I__2506 (
            .O(N__21776),
            .I(N__21773));
    LocalMux I__2505 (
            .O(N__21773),
            .I(N__21770));
    Span4Mux_v I__2504 (
            .O(N__21770),
            .I(N__21767));
    Odrv4 I__2503 (
            .O(N__21767),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__2502 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__2501 (
            .O(N__21761),
            .I(N__21758));
    Odrv12 I__2500 (
            .O(N__21758),
            .I(il_max_comp2_c));
    InMux I__2499 (
            .O(N__21755),
            .I(N__21752));
    LocalMux I__2498 (
            .O(N__21752),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__2497 (
            .O(N__21749),
            .I(N__21744));
    InMux I__2496 (
            .O(N__21748),
            .I(N__21741));
    InMux I__2495 (
            .O(N__21747),
            .I(N__21738));
    LocalMux I__2494 (
            .O(N__21744),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2493 (
            .O(N__21741),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2492 (
            .O(N__21738),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2491 (
            .O(N__21731),
            .I(N__21728));
    LocalMux I__2490 (
            .O(N__21728),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2489 (
            .O(N__21725),
            .I(N__21722));
    InMux I__2488 (
            .O(N__21722),
            .I(N__21719));
    LocalMux I__2487 (
            .O(N__21719),
            .I(N__21716));
    Odrv4 I__2486 (
            .O(N__21716),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    InMux I__2485 (
            .O(N__21713),
            .I(N__21708));
    InMux I__2484 (
            .O(N__21712),
            .I(N__21705));
    InMux I__2483 (
            .O(N__21711),
            .I(N__21702));
    LocalMux I__2482 (
            .O(N__21708),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2481 (
            .O(N__21705),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2480 (
            .O(N__21702),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2479 (
            .O(N__21695),
            .I(N__21692));
    LocalMux I__2478 (
            .O(N__21692),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2477 (
            .O(N__21689),
            .I(N__21686));
    InMux I__2476 (
            .O(N__21686),
            .I(N__21683));
    LocalMux I__2475 (
            .O(N__21683),
            .I(N__21680));
    Span4Mux_v I__2474 (
            .O(N__21680),
            .I(N__21677));
    Odrv4 I__2473 (
            .O(N__21677),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__2472 (
            .O(N__21674),
            .I(N__21669));
    InMux I__2471 (
            .O(N__21673),
            .I(N__21666));
    InMux I__2470 (
            .O(N__21672),
            .I(N__21663));
    LocalMux I__2469 (
            .O(N__21669),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2468 (
            .O(N__21666),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2467 (
            .O(N__21663),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2466 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__2465 (
            .O(N__21653),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__2464 (
            .O(N__21650),
            .I(N__21647));
    InMux I__2463 (
            .O(N__21647),
            .I(N__21644));
    LocalMux I__2462 (
            .O(N__21644),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__2461 (
            .O(N__21641),
            .I(N__21636));
    InMux I__2460 (
            .O(N__21640),
            .I(N__21633));
    InMux I__2459 (
            .O(N__21639),
            .I(N__21630));
    LocalMux I__2458 (
            .O(N__21636),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2457 (
            .O(N__21633),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2456 (
            .O(N__21630),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2455 (
            .O(N__21623),
            .I(N__21620));
    LocalMux I__2454 (
            .O(N__21620),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__2453 (
            .O(N__21617),
            .I(N__21612));
    InMux I__2452 (
            .O(N__21616),
            .I(N__21609));
    InMux I__2451 (
            .O(N__21615),
            .I(N__21606));
    LocalMux I__2450 (
            .O(N__21612),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2449 (
            .O(N__21609),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2448 (
            .O(N__21606),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__2447 (
            .O(N__21599),
            .I(N__21596));
    InMux I__2446 (
            .O(N__21596),
            .I(N__21593));
    LocalMux I__2445 (
            .O(N__21593),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2444 (
            .O(N__21590),
            .I(N__21587));
    LocalMux I__2443 (
            .O(N__21587),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2442 (
            .O(N__21584),
            .I(N__21581));
    InMux I__2441 (
            .O(N__21581),
            .I(N__21578));
    LocalMux I__2440 (
            .O(N__21578),
            .I(N__21575));
    Span4Mux_v I__2439 (
            .O(N__21575),
            .I(N__21572));
    Odrv4 I__2438 (
            .O(N__21572),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2437 (
            .O(N__21569),
            .I(N__21564));
    InMux I__2436 (
            .O(N__21568),
            .I(N__21561));
    InMux I__2435 (
            .O(N__21567),
            .I(N__21558));
    LocalMux I__2434 (
            .O(N__21564),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2433 (
            .O(N__21561),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2432 (
            .O(N__21558),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2431 (
            .O(N__21551),
            .I(N__21548));
    LocalMux I__2430 (
            .O(N__21548),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2429 (
            .O(N__21545),
            .I(N__21542));
    InMux I__2428 (
            .O(N__21542),
            .I(N__21539));
    LocalMux I__2427 (
            .O(N__21539),
            .I(N__21536));
    Span4Mux_h I__2426 (
            .O(N__21536),
            .I(N__21533));
    Odrv4 I__2425 (
            .O(N__21533),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2424 (
            .O(N__21530),
            .I(N__21525));
    InMux I__2423 (
            .O(N__21529),
            .I(N__21522));
    InMux I__2422 (
            .O(N__21528),
            .I(N__21519));
    LocalMux I__2421 (
            .O(N__21525),
            .I(N__21516));
    LocalMux I__2420 (
            .O(N__21522),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2419 (
            .O(N__21519),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2418 (
            .O(N__21516),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2417 (
            .O(N__21509),
            .I(N__21506));
    LocalMux I__2416 (
            .O(N__21506),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__2415 (
            .O(N__21503),
            .I(N__21500));
    LocalMux I__2414 (
            .O(N__21500),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2413 (
            .O(N__21497),
            .I(N__21494));
    LocalMux I__2412 (
            .O(N__21494),
            .I(N__21491));
    Odrv12 I__2411 (
            .O(N__21491),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2410 (
            .O(N__21488),
            .I(N__21485));
    LocalMux I__2409 (
            .O(N__21485),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2408 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__2407 (
            .O(N__21479),
            .I(N__21476));
    Span4Mux_v I__2406 (
            .O(N__21476),
            .I(N__21473));
    Odrv4 I__2405 (
            .O(N__21473),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2404 (
            .O(N__21470),
            .I(N__21467));
    LocalMux I__2403 (
            .O(N__21467),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__2402 (
            .O(N__21464),
            .I(N__21461));
    LocalMux I__2401 (
            .O(N__21461),
            .I(N__21458));
    Odrv4 I__2400 (
            .O(N__21458),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2399 (
            .O(N__21455),
            .I(N__21452));
    LocalMux I__2398 (
            .O(N__21452),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2397 (
            .O(N__21449),
            .I(N__21446));
    LocalMux I__2396 (
            .O(N__21446),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__2395 (
            .O(N__21443),
            .I(N__21440));
    LocalMux I__2394 (
            .O(N__21440),
            .I(N__21437));
    Odrv12 I__2393 (
            .O(N__21437),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2392 (
            .O(N__21434),
            .I(N__21431));
    LocalMux I__2391 (
            .O(N__21431),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2390 (
            .O(N__21428),
            .I(N__21425));
    LocalMux I__2389 (
            .O(N__21425),
            .I(N__21422));
    Odrv4 I__2388 (
            .O(N__21422),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    CascadeMux I__2387 (
            .O(N__21419),
            .I(N__21415));
    CascadeMux I__2386 (
            .O(N__21418),
            .I(N__21412));
    InMux I__2385 (
            .O(N__21415),
            .I(N__21399));
    InMux I__2384 (
            .O(N__21412),
            .I(N__21399));
    InMux I__2383 (
            .O(N__21411),
            .I(N__21396));
    InMux I__2382 (
            .O(N__21410),
            .I(N__21391));
    InMux I__2381 (
            .O(N__21409),
            .I(N__21391));
    InMux I__2380 (
            .O(N__21408),
            .I(N__21388));
    InMux I__2379 (
            .O(N__21407),
            .I(N__21379));
    InMux I__2378 (
            .O(N__21406),
            .I(N__21379));
    InMux I__2377 (
            .O(N__21405),
            .I(N__21379));
    InMux I__2376 (
            .O(N__21404),
            .I(N__21379));
    LocalMux I__2375 (
            .O(N__21399),
            .I(N__21372));
    LocalMux I__2374 (
            .O(N__21396),
            .I(N__21372));
    LocalMux I__2373 (
            .O(N__21391),
            .I(N__21372));
    LocalMux I__2372 (
            .O(N__21388),
            .I(N__21369));
    LocalMux I__2371 (
            .O(N__21379),
            .I(N__21364));
    Span4Mux_v I__2370 (
            .O(N__21372),
            .I(N__21364));
    Odrv4 I__2369 (
            .O(N__21369),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2368 (
            .O(N__21364),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2367 (
            .O(N__21359),
            .I(N__21352));
    CascadeMux I__2366 (
            .O(N__21358),
            .I(N__21349));
    InMux I__2365 (
            .O(N__21357),
            .I(N__21343));
    InMux I__2364 (
            .O(N__21356),
            .I(N__21334));
    InMux I__2363 (
            .O(N__21355),
            .I(N__21334));
    InMux I__2362 (
            .O(N__21352),
            .I(N__21334));
    InMux I__2361 (
            .O(N__21349),
            .I(N__21334));
    CascadeMux I__2360 (
            .O(N__21348),
            .I(N__21331));
    CascadeMux I__2359 (
            .O(N__21347),
            .I(N__21327));
    CascadeMux I__2358 (
            .O(N__21346),
            .I(N__21324));
    LocalMux I__2357 (
            .O(N__21343),
            .I(N__21318));
    LocalMux I__2356 (
            .O(N__21334),
            .I(N__21318));
    InMux I__2355 (
            .O(N__21331),
            .I(N__21311));
    InMux I__2354 (
            .O(N__21330),
            .I(N__21311));
    InMux I__2353 (
            .O(N__21327),
            .I(N__21311));
    InMux I__2352 (
            .O(N__21324),
            .I(N__21308));
    InMux I__2351 (
            .O(N__21323),
            .I(N__21305));
    Span4Mux_v I__2350 (
            .O(N__21318),
            .I(N__21298));
    LocalMux I__2349 (
            .O(N__21311),
            .I(N__21298));
    LocalMux I__2348 (
            .O(N__21308),
            .I(N__21298));
    LocalMux I__2347 (
            .O(N__21305),
            .I(N__21295));
    Odrv4 I__2346 (
            .O(N__21298),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2345 (
            .O(N__21295),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__2344 (
            .O(N__21290),
            .I(N__21283));
    InMux I__2343 (
            .O(N__21289),
            .I(N__21274));
    InMux I__2342 (
            .O(N__21288),
            .I(N__21274));
    InMux I__2341 (
            .O(N__21287),
            .I(N__21274));
    InMux I__2340 (
            .O(N__21286),
            .I(N__21274));
    InMux I__2339 (
            .O(N__21283),
            .I(N__21270));
    LocalMux I__2338 (
            .O(N__21274),
            .I(N__21266));
    CascadeMux I__2337 (
            .O(N__21273),
            .I(N__21258));
    LocalMux I__2336 (
            .O(N__21270),
            .I(N__21255));
    CascadeMux I__2335 (
            .O(N__21269),
            .I(N__21241));
    Span4Mux_h I__2334 (
            .O(N__21266),
            .I(N__21238));
    InMux I__2333 (
            .O(N__21265),
            .I(N__21233));
    InMux I__2332 (
            .O(N__21264),
            .I(N__21233));
    InMux I__2331 (
            .O(N__21263),
            .I(N__21226));
    InMux I__2330 (
            .O(N__21262),
            .I(N__21226));
    InMux I__2329 (
            .O(N__21261),
            .I(N__21226));
    InMux I__2328 (
            .O(N__21258),
            .I(N__21223));
    Span4Mux_v I__2327 (
            .O(N__21255),
            .I(N__21220));
    InMux I__2326 (
            .O(N__21254),
            .I(N__21213));
    InMux I__2325 (
            .O(N__21253),
            .I(N__21213));
    InMux I__2324 (
            .O(N__21252),
            .I(N__21213));
    InMux I__2323 (
            .O(N__21251),
            .I(N__21196));
    InMux I__2322 (
            .O(N__21250),
            .I(N__21196));
    InMux I__2321 (
            .O(N__21249),
            .I(N__21196));
    InMux I__2320 (
            .O(N__21248),
            .I(N__21196));
    InMux I__2319 (
            .O(N__21247),
            .I(N__21196));
    InMux I__2318 (
            .O(N__21246),
            .I(N__21196));
    InMux I__2317 (
            .O(N__21245),
            .I(N__21196));
    InMux I__2316 (
            .O(N__21244),
            .I(N__21196));
    InMux I__2315 (
            .O(N__21241),
            .I(N__21193));
    Span4Mux_v I__2314 (
            .O(N__21238),
            .I(N__21186));
    LocalMux I__2313 (
            .O(N__21233),
            .I(N__21186));
    LocalMux I__2312 (
            .O(N__21226),
            .I(N__21186));
    LocalMux I__2311 (
            .O(N__21223),
            .I(N__21179));
    Sp12to4 I__2310 (
            .O(N__21220),
            .I(N__21179));
    LocalMux I__2309 (
            .O(N__21213),
            .I(N__21179));
    LocalMux I__2308 (
            .O(N__21196),
            .I(N__21167));
    LocalMux I__2307 (
            .O(N__21193),
            .I(N__21164));
    Span4Mux_s2_h I__2306 (
            .O(N__21186),
            .I(N__21161));
    Span12Mux_h I__2305 (
            .O(N__21179),
            .I(N__21158));
    InMux I__2304 (
            .O(N__21178),
            .I(N__21155));
    InMux I__2303 (
            .O(N__21177),
            .I(N__21152));
    InMux I__2302 (
            .O(N__21176),
            .I(N__21137));
    InMux I__2301 (
            .O(N__21175),
            .I(N__21137));
    InMux I__2300 (
            .O(N__21174),
            .I(N__21137));
    InMux I__2299 (
            .O(N__21173),
            .I(N__21137));
    InMux I__2298 (
            .O(N__21172),
            .I(N__21137));
    InMux I__2297 (
            .O(N__21171),
            .I(N__21137));
    InMux I__2296 (
            .O(N__21170),
            .I(N__21137));
    Span4Mux_s1_h I__2295 (
            .O(N__21167),
            .I(N__21134));
    Span4Mux_v I__2294 (
            .O(N__21164),
            .I(N__21129));
    Span4Mux_v I__2293 (
            .O(N__21161),
            .I(N__21129));
    Odrv12 I__2292 (
            .O(N__21158),
            .I(N_19_1));
    LocalMux I__2291 (
            .O(N__21155),
            .I(N_19_1));
    LocalMux I__2290 (
            .O(N__21152),
            .I(N_19_1));
    LocalMux I__2289 (
            .O(N__21137),
            .I(N_19_1));
    Odrv4 I__2288 (
            .O(N__21134),
            .I(N_19_1));
    Odrv4 I__2287 (
            .O(N__21129),
            .I(N_19_1));
    InMux I__2286 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__2285 (
            .O(N__21113),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    CascadeMux I__2284 (
            .O(N__21110),
            .I(N__21107));
    InMux I__2283 (
            .O(N__21107),
            .I(N__21104));
    LocalMux I__2282 (
            .O(N__21104),
            .I(N__21101));
    Span4Mux_h I__2281 (
            .O(N__21101),
            .I(N__21098));
    Odrv4 I__2280 (
            .O(N__21098),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__2279 (
            .O(N__21095),
            .I(N__21090));
    InMux I__2278 (
            .O(N__21094),
            .I(N__21087));
    InMux I__2277 (
            .O(N__21093),
            .I(N__21084));
    LocalMux I__2276 (
            .O(N__21090),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2275 (
            .O(N__21087),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2274 (
            .O(N__21084),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2273 (
            .O(N__21077),
            .I(N__21074));
    LocalMux I__2272 (
            .O(N__21074),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__2271 (
            .O(N__21071),
            .I(N__21066));
    InMux I__2270 (
            .O(N__21070),
            .I(N__21063));
    InMux I__2269 (
            .O(N__21069),
            .I(N__21060));
    LocalMux I__2268 (
            .O(N__21066),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2267 (
            .O(N__21063),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2266 (
            .O(N__21060),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__2265 (
            .O(N__21053),
            .I(N__21050));
    InMux I__2264 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__2263 (
            .O(N__21047),
            .I(N__21044));
    Span4Mux_s3_h I__2262 (
            .O(N__21044),
            .I(N__21041));
    Odrv4 I__2261 (
            .O(N__21041),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2260 (
            .O(N__21038),
            .I(N__21034));
    InMux I__2259 (
            .O(N__21037),
            .I(N__21030));
    LocalMux I__2258 (
            .O(N__21034),
            .I(N__21027));
    InMux I__2257 (
            .O(N__21033),
            .I(N__21024));
    LocalMux I__2256 (
            .O(N__21030),
            .I(N__21017));
    Span4Mux_h I__2255 (
            .O(N__21027),
            .I(N__21017));
    LocalMux I__2254 (
            .O(N__21024),
            .I(N__21017));
    Odrv4 I__2253 (
            .O(N__21017),
            .I(pwm_duty_input_7));
    InMux I__2252 (
            .O(N__21014),
            .I(N__21011));
    LocalMux I__2251 (
            .O(N__21011),
            .I(N__21007));
    InMux I__2250 (
            .O(N__21010),
            .I(N__21003));
    Span4Mux_h I__2249 (
            .O(N__21007),
            .I(N__21000));
    InMux I__2248 (
            .O(N__21006),
            .I(N__20997));
    LocalMux I__2247 (
            .O(N__21003),
            .I(pwm_duty_input_5));
    Odrv4 I__2246 (
            .O(N__21000),
            .I(pwm_duty_input_5));
    LocalMux I__2245 (
            .O(N__20997),
            .I(pwm_duty_input_5));
    CascadeMux I__2244 (
            .O(N__20990),
            .I(N__20987));
    InMux I__2243 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__2242 (
            .O(N__20984),
            .I(N__20981));
    Odrv12 I__2241 (
            .O(N__20981),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ));
    InMux I__2240 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__2239 (
            .O(N__20975),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2238 (
            .O(N__20972),
            .I(N__20969));
    LocalMux I__2237 (
            .O(N__20969),
            .I(N__20966));
    Odrv4 I__2236 (
            .O(N__20966),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2235 (
            .O(N__20963),
            .I(N__20960));
    LocalMux I__2234 (
            .O(N__20960),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2233 (
            .O(N__20957),
            .I(N__20954));
    LocalMux I__2232 (
            .O(N__20954),
            .I(N__20951));
    Odrv4 I__2231 (
            .O(N__20951),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2230 (
            .O(N__20948),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2229 (
            .O(N__20945),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2228 (
            .O(N__20942),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2227 (
            .O(N__20939),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2226 (
            .O(N__20936),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2225 (
            .O(N__20933),
            .I(bfn_3_10_0_));
    InMux I__2224 (
            .O(N__20930),
            .I(N__20916));
    InMux I__2223 (
            .O(N__20929),
            .I(N__20916));
    InMux I__2222 (
            .O(N__20928),
            .I(N__20916));
    InMux I__2221 (
            .O(N__20927),
            .I(N__20916));
    InMux I__2220 (
            .O(N__20926),
            .I(N__20909));
    InMux I__2219 (
            .O(N__20925),
            .I(N__20906));
    LocalMux I__2218 (
            .O(N__20916),
            .I(N__20903));
    InMux I__2217 (
            .O(N__20915),
            .I(N__20894));
    InMux I__2216 (
            .O(N__20914),
            .I(N__20894));
    InMux I__2215 (
            .O(N__20913),
            .I(N__20894));
    InMux I__2214 (
            .O(N__20912),
            .I(N__20894));
    LocalMux I__2213 (
            .O(N__20909),
            .I(N__20889));
    LocalMux I__2212 (
            .O(N__20906),
            .I(N__20889));
    Odrv4 I__2211 (
            .O(N__20903),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2210 (
            .O(N__20894),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__2209 (
            .O(N__20889),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2208 (
            .O(N__20882),
            .I(\pwm_generator_inst.counter_cry_8 ));
    CascadeMux I__2207 (
            .O(N__20879),
            .I(N__20876));
    InMux I__2206 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2205 (
            .O(N__20873),
            .I(N__20869));
    InMux I__2204 (
            .O(N__20872),
            .I(N__20866));
    Span4Mux_s2_h I__2203 (
            .O(N__20869),
            .I(N__20863));
    LocalMux I__2202 (
            .O(N__20866),
            .I(N__20860));
    Odrv4 I__2201 (
            .O(N__20863),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    Odrv12 I__2200 (
            .O(N__20860),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__2199 (
            .O(N__20855),
            .I(N__20850));
    CascadeMux I__2198 (
            .O(N__20854),
            .I(N__20847));
    InMux I__2197 (
            .O(N__20853),
            .I(N__20844));
    LocalMux I__2196 (
            .O(N__20850),
            .I(N__20841));
    InMux I__2195 (
            .O(N__20847),
            .I(N__20838));
    LocalMux I__2194 (
            .O(N__20844),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    Odrv4 I__2193 (
            .O(N__20841),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2192 (
            .O(N__20838),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    CascadeMux I__2191 (
            .O(N__20831),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__2190 (
            .O(N__20828),
            .I(N__20825));
    LocalMux I__2189 (
            .O(N__20825),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__2188 (
            .O(N__20822),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__2187 (
            .O(N__20819),
            .I(bfn_3_9_0_));
    InMux I__2186 (
            .O(N__20816),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2185 (
            .O(N__20813),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2184 (
            .O(N__20810),
            .I(N__20807));
    LocalMux I__2183 (
            .O(N__20807),
            .I(N__20804));
    Span4Mux_h I__2182 (
            .O(N__20804),
            .I(N__20801));
    Span4Mux_v I__2181 (
            .O(N__20801),
            .I(N__20798));
    Odrv4 I__2180 (
            .O(N__20798),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2179 (
            .O(N__20795),
            .I(bfn_2_17_0_));
    InMux I__2178 (
            .O(N__20792),
            .I(N__20789));
    LocalMux I__2177 (
            .O(N__20789),
            .I(N__20786));
    Odrv4 I__2176 (
            .O(N__20786),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    CascadeMux I__2175 (
            .O(N__20783),
            .I(N__20780));
    InMux I__2174 (
            .O(N__20780),
            .I(N__20777));
    LocalMux I__2173 (
            .O(N__20777),
            .I(N__20774));
    Odrv12 I__2172 (
            .O(N__20774),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2171 (
            .O(N__20771),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    InMux I__2170 (
            .O(N__20768),
            .I(N__20764));
    InMux I__2169 (
            .O(N__20767),
            .I(N__20761));
    LocalMux I__2168 (
            .O(N__20764),
            .I(N__20758));
    LocalMux I__2167 (
            .O(N__20761),
            .I(N__20755));
    Odrv4 I__2166 (
            .O(N__20758),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    Odrv12 I__2165 (
            .O(N__20755),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    InMux I__2164 (
            .O(N__20750),
            .I(N__20745));
    InMux I__2163 (
            .O(N__20749),
            .I(N__20742));
    InMux I__2162 (
            .O(N__20748),
            .I(N__20739));
    LocalMux I__2161 (
            .O(N__20745),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__2160 (
            .O(N__20742),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__2159 (
            .O(N__20739),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__2158 (
            .O(N__20732),
            .I(N__20728));
    InMux I__2157 (
            .O(N__20731),
            .I(N__20725));
    LocalMux I__2156 (
            .O(N__20728),
            .I(N__20722));
    LocalMux I__2155 (
            .O(N__20725),
            .I(N__20719));
    Odrv4 I__2154 (
            .O(N__20722),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    Odrv12 I__2153 (
            .O(N__20719),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    InMux I__2152 (
            .O(N__20714),
            .I(N__20709));
    InMux I__2151 (
            .O(N__20713),
            .I(N__20706));
    InMux I__2150 (
            .O(N__20712),
            .I(N__20703));
    LocalMux I__2149 (
            .O(N__20709),
            .I(N__20700));
    LocalMux I__2148 (
            .O(N__20706),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2147 (
            .O(N__20703),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    Odrv4 I__2146 (
            .O(N__20700),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__2145 (
            .O(N__20693),
            .I(N__20689));
    InMux I__2144 (
            .O(N__20692),
            .I(N__20686));
    LocalMux I__2143 (
            .O(N__20689),
            .I(N__20683));
    LocalMux I__2142 (
            .O(N__20686),
            .I(N__20680));
    Odrv4 I__2141 (
            .O(N__20683),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    Odrv12 I__2140 (
            .O(N__20680),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__2139 (
            .O(N__20675),
            .I(N__20672));
    LocalMux I__2138 (
            .O(N__20672),
            .I(N__20668));
    InMux I__2137 (
            .O(N__20671),
            .I(N__20664));
    Span4Mux_s2_h I__2136 (
            .O(N__20668),
            .I(N__20661));
    InMux I__2135 (
            .O(N__20667),
            .I(N__20658));
    LocalMux I__2134 (
            .O(N__20664),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__2133 (
            .O(N__20661),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2132 (
            .O(N__20658),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__2131 (
            .O(N__20651),
            .I(N__20647));
    InMux I__2130 (
            .O(N__20650),
            .I(N__20644));
    LocalMux I__2129 (
            .O(N__20647),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__2128 (
            .O(N__20644),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2127 (
            .O(N__20639),
            .I(N__20633));
    InMux I__2126 (
            .O(N__20638),
            .I(N__20633));
    LocalMux I__2125 (
            .O(N__20633),
            .I(N__20630));
    Odrv12 I__2124 (
            .O(N__20630),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    InMux I__2123 (
            .O(N__20627),
            .I(N__20624));
    LocalMux I__2122 (
            .O(N__20624),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    CascadeMux I__2121 (
            .O(N__20621),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ));
    InMux I__2120 (
            .O(N__20618),
            .I(N__20613));
    CascadeMux I__2119 (
            .O(N__20617),
            .I(N__20608));
    InMux I__2118 (
            .O(N__20616),
            .I(N__20605));
    LocalMux I__2117 (
            .O(N__20613),
            .I(N__20602));
    InMux I__2116 (
            .O(N__20612),
            .I(N__20593));
    InMux I__2115 (
            .O(N__20611),
            .I(N__20590));
    InMux I__2114 (
            .O(N__20608),
            .I(N__20587));
    LocalMux I__2113 (
            .O(N__20605),
            .I(N__20582));
    Span4Mux_v I__2112 (
            .O(N__20602),
            .I(N__20582));
    InMux I__2111 (
            .O(N__20601),
            .I(N__20579));
    InMux I__2110 (
            .O(N__20600),
            .I(N__20568));
    InMux I__2109 (
            .O(N__20599),
            .I(N__20568));
    InMux I__2108 (
            .O(N__20598),
            .I(N__20568));
    InMux I__2107 (
            .O(N__20597),
            .I(N__20568));
    InMux I__2106 (
            .O(N__20596),
            .I(N__20568));
    LocalMux I__2105 (
            .O(N__20593),
            .I(N__20565));
    LocalMux I__2104 (
            .O(N__20590),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2103 (
            .O(N__20587),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2102 (
            .O(N__20582),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2101 (
            .O(N__20579),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2100 (
            .O(N__20568),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv12 I__2099 (
            .O(N__20565),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    CascadeMux I__2098 (
            .O(N__20552),
            .I(N__20549));
    InMux I__2097 (
            .O(N__20549),
            .I(N__20546));
    LocalMux I__2096 (
            .O(N__20546),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__2095 (
            .O(N__20543),
            .I(N__20540));
    LocalMux I__2094 (
            .O(N__20540),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    InMux I__2093 (
            .O(N__20537),
            .I(N__20534));
    LocalMux I__2092 (
            .O(N__20534),
            .I(N__20531));
    Odrv4 I__2091 (
            .O(N__20531),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2090 (
            .O(N__20528),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__2089 (
            .O(N__20525),
            .I(N__20522));
    LocalMux I__2088 (
            .O(N__20522),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__2087 (
            .O(N__20519),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    CascadeMux I__2086 (
            .O(N__20516),
            .I(N__20513));
    InMux I__2085 (
            .O(N__20513),
            .I(N__20510));
    LocalMux I__2084 (
            .O(N__20510),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__2083 (
            .O(N__20507),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__2082 (
            .O(N__20504),
            .I(N__20501));
    LocalMux I__2081 (
            .O(N__20501),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__2080 (
            .O(N__20498),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__2079 (
            .O(N__20495),
            .I(N__20492));
    LocalMux I__2078 (
            .O(N__20492),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__2077 (
            .O(N__20489),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__2076 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__2075 (
            .O(N__20483),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__2074 (
            .O(N__20480),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__2073 (
            .O(N__20477),
            .I(N__20474));
    LocalMux I__2072 (
            .O(N__20474),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2071 (
            .O(N__20471),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__2070 (
            .O(N__20468),
            .I(N__20465));
    LocalMux I__2069 (
            .O(N__20465),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__2068 (
            .O(N__20462),
            .I(N__20459));
    LocalMux I__2067 (
            .O(N__20459),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__2066 (
            .O(N__20456),
            .I(N__20453));
    LocalMux I__2065 (
            .O(N__20453),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__2064 (
            .O(N__20450),
            .I(N__20447));
    LocalMux I__2063 (
            .O(N__20447),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__2062 (
            .O(N__20444),
            .I(N__20441));
    LocalMux I__2061 (
            .O(N__20441),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__2060 (
            .O(N__20438),
            .I(N__20435));
    LocalMux I__2059 (
            .O(N__20435),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__2058 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__2057 (
            .O(N__20429),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__2056 (
            .O(N__20426),
            .I(N__20423));
    LocalMux I__2055 (
            .O(N__20423),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__2054 (
            .O(N__20420),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    CascadeMux I__2053 (
            .O(N__20417),
            .I(N__20414));
    InMux I__2052 (
            .O(N__20414),
            .I(N__20411));
    LocalMux I__2051 (
            .O(N__20411),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__2050 (
            .O(N__20408),
            .I(N__20405));
    LocalMux I__2049 (
            .O(N__20405),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__2048 (
            .O(N__20402),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    CascadeMux I__2047 (
            .O(N__20399),
            .I(N__20396));
    InMux I__2046 (
            .O(N__20396),
            .I(N__20393));
    LocalMux I__2045 (
            .O(N__20393),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__2044 (
            .O(N__20390),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__2043 (
            .O(N__20387),
            .I(N__20384));
    LocalMux I__2042 (
            .O(N__20384),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__2041 (
            .O(N__20381),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__2040 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__2039 (
            .O(N__20375),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__2038 (
            .O(N__20372),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__2037 (
            .O(N__20369),
            .I(N__20366));
    LocalMux I__2036 (
            .O(N__20366),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__2035 (
            .O(N__20363),
            .I(bfn_2_14_0_));
    InMux I__2034 (
            .O(N__20360),
            .I(N__20357));
    LocalMux I__2033 (
            .O(N__20357),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__2032 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__2031 (
            .O(N__20351),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__2030 (
            .O(N__20348),
            .I(N__20345));
    LocalMux I__2029 (
            .O(N__20345),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    CascadeMux I__2028 (
            .O(N__20342),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__2027 (
            .O(N__20339),
            .I(N__20334));
    InMux I__2026 (
            .O(N__20338),
            .I(N__20329));
    InMux I__2025 (
            .O(N__20337),
            .I(N__20329));
    LocalMux I__2024 (
            .O(N__20334),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2023 (
            .O(N__20329),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__2022 (
            .O(N__20324),
            .I(N__20320));
    InMux I__2021 (
            .O(N__20323),
            .I(N__20316));
    InMux I__2020 (
            .O(N__20320),
            .I(N__20313));
    InMux I__2019 (
            .O(N__20319),
            .I(N__20310));
    LocalMux I__2018 (
            .O(N__20316),
            .I(N__20307));
    LocalMux I__2017 (
            .O(N__20313),
            .I(N__20302));
    LocalMux I__2016 (
            .O(N__20310),
            .I(N__20302));
    Odrv4 I__2015 (
            .O(N__20307),
            .I(pwm_duty_input_9));
    Odrv4 I__2014 (
            .O(N__20302),
            .I(pwm_duty_input_9));
    InMux I__2013 (
            .O(N__20297),
            .I(N__20292));
    InMux I__2012 (
            .O(N__20296),
            .I(N__20289));
    InMux I__2011 (
            .O(N__20295),
            .I(N__20286));
    LocalMux I__2010 (
            .O(N__20292),
            .I(pwm_duty_input_6));
    LocalMux I__2009 (
            .O(N__20289),
            .I(pwm_duty_input_6));
    LocalMux I__2008 (
            .O(N__20286),
            .I(pwm_duty_input_6));
    InMux I__2007 (
            .O(N__20279),
            .I(N__20276));
    LocalMux I__2006 (
            .O(N__20276),
            .I(N__20273));
    Odrv4 I__2005 (
            .O(N__20273),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    CascadeMux I__2004 (
            .O(N__20270),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ));
    InMux I__2003 (
            .O(N__20267),
            .I(N__20262));
    InMux I__2002 (
            .O(N__20266),
            .I(N__20259));
    InMux I__2001 (
            .O(N__20265),
            .I(N__20256));
    LocalMux I__2000 (
            .O(N__20262),
            .I(pwm_duty_input_8));
    LocalMux I__1999 (
            .O(N__20259),
            .I(pwm_duty_input_8));
    LocalMux I__1998 (
            .O(N__20256),
            .I(pwm_duty_input_8));
    InMux I__1997 (
            .O(N__20249),
            .I(N__20244));
    InMux I__1996 (
            .O(N__20248),
            .I(N__20239));
    InMux I__1995 (
            .O(N__20247),
            .I(N__20239));
    LocalMux I__1994 (
            .O(N__20244),
            .I(N__20236));
    LocalMux I__1993 (
            .O(N__20239),
            .I(N__20233));
    Span4Mux_s1_h I__1992 (
            .O(N__20236),
            .I(N__20230));
    Odrv4 I__1991 (
            .O(N__20233),
            .I(pwm_duty_input_3));
    Odrv4 I__1990 (
            .O(N__20230),
            .I(pwm_duty_input_3));
    CascadeMux I__1989 (
            .O(N__20225),
            .I(N__20222));
    InMux I__1988 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__1987 (
            .O(N__20219),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__1986 (
            .O(N__20216),
            .I(N__20210));
    InMux I__1985 (
            .O(N__20215),
            .I(N__20210));
    LocalMux I__1984 (
            .O(N__20210),
            .I(N__20206));
    InMux I__1983 (
            .O(N__20209),
            .I(N__20203));
    Span4Mux_h I__1982 (
            .O(N__20206),
            .I(N__20198));
    LocalMux I__1981 (
            .O(N__20203),
            .I(N__20198));
    Span4Mux_s1_h I__1980 (
            .O(N__20198),
            .I(N__20195));
    Odrv4 I__1979 (
            .O(N__20195),
            .I(pwm_duty_input_4));
    InMux I__1978 (
            .O(N__20192),
            .I(N__20188));
    InMux I__1977 (
            .O(N__20191),
            .I(N__20185));
    LocalMux I__1976 (
            .O(N__20188),
            .I(N__20182));
    LocalMux I__1975 (
            .O(N__20185),
            .I(N__20179));
    Span4Mux_v I__1974 (
            .O(N__20182),
            .I(N__20176));
    Span4Mux_v I__1973 (
            .O(N__20179),
            .I(N__20173));
    Odrv4 I__1972 (
            .O(N__20176),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    Odrv4 I__1971 (
            .O(N__20173),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1970 (
            .O(N__20168),
            .I(N__20165));
    LocalMux I__1969 (
            .O(N__20165),
            .I(N__20162));
    Span4Mux_h I__1968 (
            .O(N__20162),
            .I(N__20159));
    Odrv4 I__1967 (
            .O(N__20159),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1966 (
            .O(N__20156),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1965 (
            .O(N__20153),
            .I(N__20150));
    LocalMux I__1964 (
            .O(N__20150),
            .I(N__20147));
    Span4Mux_h I__1963 (
            .O(N__20147),
            .I(N__20144));
    Odrv4 I__1962 (
            .O(N__20144),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1961 (
            .O(N__20141),
            .I(N__20138));
    LocalMux I__1960 (
            .O(N__20138),
            .I(N__20135));
    Span4Mux_v I__1959 (
            .O(N__20135),
            .I(N__20131));
    InMux I__1958 (
            .O(N__20134),
            .I(N__20128));
    Odrv4 I__1957 (
            .O(N__20131),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    LocalMux I__1956 (
            .O(N__20128),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__1955 (
            .O(N__20123),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1954 (
            .O(N__20120),
            .I(N__20117));
    LocalMux I__1953 (
            .O(N__20117),
            .I(N__20114));
    Span4Mux_h I__1952 (
            .O(N__20114),
            .I(N__20111));
    Odrv4 I__1951 (
            .O(N__20111),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1950 (
            .O(N__20108),
            .I(N__20105));
    LocalMux I__1949 (
            .O(N__20105),
            .I(N__20101));
    InMux I__1948 (
            .O(N__20104),
            .I(N__20098));
    Span4Mux_s2_h I__1947 (
            .O(N__20101),
            .I(N__20093));
    LocalMux I__1946 (
            .O(N__20098),
            .I(N__20093));
    Odrv4 I__1945 (
            .O(N__20093),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__1944 (
            .O(N__20090),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    CascadeMux I__1943 (
            .O(N__20087),
            .I(\current_shift_inst.PI_CTRL.N_168_cascade_ ));
    CascadeMux I__1942 (
            .O(N__20084),
            .I(N__20079));
    CascadeMux I__1941 (
            .O(N__20083),
            .I(N__20076));
    InMux I__1940 (
            .O(N__20082),
            .I(N__20066));
    InMux I__1939 (
            .O(N__20079),
            .I(N__20066));
    InMux I__1938 (
            .O(N__20076),
            .I(N__20066));
    InMux I__1937 (
            .O(N__20075),
            .I(N__20066));
    LocalMux I__1936 (
            .O(N__20066),
            .I(\current_shift_inst.PI_CTRL.N_166 ));
    InMux I__1935 (
            .O(N__20063),
            .I(N__20059));
    InMux I__1934 (
            .O(N__20062),
            .I(N__20055));
    LocalMux I__1933 (
            .O(N__20059),
            .I(N__20052));
    InMux I__1932 (
            .O(N__20058),
            .I(N__20049));
    LocalMux I__1931 (
            .O(N__20055),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__1930 (
            .O(N__20052),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    LocalMux I__1929 (
            .O(N__20049),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__1928 (
            .O(N__20042),
            .I(N__20039));
    LocalMux I__1927 (
            .O(N__20039),
            .I(N__20035));
    InMux I__1926 (
            .O(N__20038),
            .I(N__20032));
    Odrv4 I__1925 (
            .O(N__20035),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    LocalMux I__1924 (
            .O(N__20032),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1923 (
            .O(N__20027),
            .I(\current_shift_inst.PI_CTRL.N_166_cascade_ ));
    InMux I__1922 (
            .O(N__20024),
            .I(N__20015));
    InMux I__1921 (
            .O(N__20023),
            .I(N__20015));
    InMux I__1920 (
            .O(N__20022),
            .I(N__20015));
    LocalMux I__1919 (
            .O(N__20015),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1918 (
            .O(N__20012),
            .I(N__20009));
    LocalMux I__1917 (
            .O(N__20009),
            .I(\current_shift_inst.PI_CTRL.N_162 ));
    InMux I__1916 (
            .O(N__20006),
            .I(N__20002));
    InMux I__1915 (
            .O(N__20005),
            .I(N__19999));
    LocalMux I__1914 (
            .O(N__20002),
            .I(N__19996));
    LocalMux I__1913 (
            .O(N__19999),
            .I(pwm_duty_input_0));
    Odrv4 I__1912 (
            .O(N__19996),
            .I(pwm_duty_input_0));
    InMux I__1911 (
            .O(N__19991),
            .I(N__19987));
    InMux I__1910 (
            .O(N__19990),
            .I(N__19984));
    LocalMux I__1909 (
            .O(N__19987),
            .I(N__19981));
    LocalMux I__1908 (
            .O(N__19984),
            .I(pwm_duty_input_1));
    Odrv4 I__1907 (
            .O(N__19981),
            .I(pwm_duty_input_1));
    InMux I__1906 (
            .O(N__19976),
            .I(N__19972));
    InMux I__1905 (
            .O(N__19975),
            .I(N__19969));
    LocalMux I__1904 (
            .O(N__19972),
            .I(N__19966));
    LocalMux I__1903 (
            .O(N__19969),
            .I(pwm_duty_input_2));
    Odrv4 I__1902 (
            .O(N__19966),
            .I(pwm_duty_input_2));
    InMux I__1901 (
            .O(N__19961),
            .I(N__19952));
    InMux I__1900 (
            .O(N__19960),
            .I(N__19952));
    InMux I__1899 (
            .O(N__19959),
            .I(N__19952));
    LocalMux I__1898 (
            .O(N__19952),
            .I(\current_shift_inst.PI_CTRL.N_167 ));
    CascadeMux I__1897 (
            .O(N__19949),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    InMux I__1896 (
            .O(N__19946),
            .I(N__19942));
    InMux I__1895 (
            .O(N__19945),
            .I(N__19939));
    LocalMux I__1894 (
            .O(N__19942),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__1893 (
            .O(N__19939),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__1892 (
            .O(N__19934),
            .I(N__19931));
    LocalMux I__1891 (
            .O(N__19931),
            .I(N__19928));
    Odrv4 I__1890 (
            .O(N__19928),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__1889 (
            .O(N__19925),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__1888 (
            .O(N__19922),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__1887 (
            .O(N__19919),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__1886 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__1885 (
            .O(N__19913),
            .I(N_34_i_i));
    InMux I__1884 (
            .O(N__19910),
            .I(N__19907));
    LocalMux I__1883 (
            .O(N__19907),
            .I(rgb_drv_RNOZ0));
    InMux I__1882 (
            .O(N__19904),
            .I(N__19901));
    LocalMux I__1881 (
            .O(N__19901),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__1880 (
            .O(N__19898),
            .I(N__19895));
    LocalMux I__1879 (
            .O(N__19895),
            .I(N__19892));
    Span4Mux_v I__1878 (
            .O(N__19892),
            .I(N__19889));
    Span4Mux_v I__1877 (
            .O(N__19889),
            .I(N__19886));
    Odrv4 I__1876 (
            .O(N__19886),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1875 (
            .O(N__19883),
            .I(N__19880));
    LocalMux I__1874 (
            .O(N__19880),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1873 (
            .O(N__19877),
            .I(N__19874));
    LocalMux I__1872 (
            .O(N__19874),
            .I(N__19870));
    InMux I__1871 (
            .O(N__19873),
            .I(N__19867));
    Span4Mux_s2_h I__1870 (
            .O(N__19870),
            .I(N__19864));
    LocalMux I__1869 (
            .O(N__19867),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__1868 (
            .O(N__19864),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    InMux I__1867 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__1866 (
            .O(N__19856),
            .I(N__19853));
    Span4Mux_v I__1865 (
            .O(N__19853),
            .I(N__19850));
    Odrv4 I__1864 (
            .O(N__19850),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__1863 (
            .O(N__19847),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1862 (
            .O(N__19844),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1861 (
            .O(N__19841),
            .I(N__19838));
    LocalMux I__1860 (
            .O(N__19838),
            .I(N__19835));
    Span4Mux_v I__1859 (
            .O(N__19835),
            .I(N__19832));
    Odrv4 I__1858 (
            .O(N__19832),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__1857 (
            .O(N__19829),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1856 (
            .O(N__19826),
            .I(N__19822));
    InMux I__1855 (
            .O(N__19825),
            .I(N__19818));
    LocalMux I__1854 (
            .O(N__19822),
            .I(N__19815));
    InMux I__1853 (
            .O(N__19821),
            .I(N__19812));
    LocalMux I__1852 (
            .O(N__19818),
            .I(N__19807));
    Span4Mux_v I__1851 (
            .O(N__19815),
            .I(N__19807));
    LocalMux I__1850 (
            .O(N__19812),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__1849 (
            .O(N__19807),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    CascadeMux I__1848 (
            .O(N__19802),
            .I(N__19799));
    InMux I__1847 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__1846 (
            .O(N__19796),
            .I(N__19793));
    Odrv4 I__1845 (
            .O(N__19793),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__1844 (
            .O(N__19790),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1843 (
            .O(N__19787),
            .I(N__19782));
    InMux I__1842 (
            .O(N__19786),
            .I(N__19779));
    InMux I__1841 (
            .O(N__19785),
            .I(N__19776));
    LocalMux I__1840 (
            .O(N__19782),
            .I(N__19773));
    LocalMux I__1839 (
            .O(N__19779),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__1838 (
            .O(N__19776),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    Odrv4 I__1837 (
            .O(N__19773),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    CascadeMux I__1836 (
            .O(N__19766),
            .I(N__19763));
    InMux I__1835 (
            .O(N__19763),
            .I(N__19760));
    LocalMux I__1834 (
            .O(N__19760),
            .I(N__19757));
    Odrv12 I__1833 (
            .O(N__19757),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__1832 (
            .O(N__19754),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    CascadeMux I__1831 (
            .O(N__19751),
            .I(N__19748));
    InMux I__1830 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__1829 (
            .O(N__19745),
            .I(N__19742));
    Odrv12 I__1828 (
            .O(N__19742),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__1827 (
            .O(N__19739),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    CascadeMux I__1826 (
            .O(N__19736),
            .I(N__19733));
    InMux I__1825 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__1824 (
            .O(N__19730),
            .I(N__19727));
    Odrv4 I__1823 (
            .O(N__19727),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__1822 (
            .O(N__19724),
            .I(bfn_1_19_0_));
    InMux I__1821 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__1820 (
            .O(N__19718),
            .I(N__19715));
    Span4Mux_v I__1819 (
            .O(N__19715),
            .I(N__19712));
    Span4Mux_v I__1818 (
            .O(N__19712),
            .I(N__19709));
    Odrv4 I__1817 (
            .O(N__19709),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1816 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__1815 (
            .O(N__19703),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1814 (
            .O(N__19700),
            .I(N__19697));
    LocalMux I__1813 (
            .O(N__19697),
            .I(N__19694));
    Span4Mux_v I__1812 (
            .O(N__19694),
            .I(N__19691));
    Odrv4 I__1811 (
            .O(N__19691),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1810 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__1809 (
            .O(N__19685),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1808 (
            .O(N__19682),
            .I(N__19679));
    LocalMux I__1807 (
            .O(N__19679),
            .I(N__19676));
    Span4Mux_h I__1806 (
            .O(N__19676),
            .I(N__19673));
    Span4Mux_v I__1805 (
            .O(N__19673),
            .I(N__19670));
    Odrv4 I__1804 (
            .O(N__19670),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1803 (
            .O(N__19667),
            .I(N__19664));
    LocalMux I__1802 (
            .O(N__19664),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1801 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__1800 (
            .O(N__19658),
            .I(N__19655));
    Span4Mux_h I__1799 (
            .O(N__19655),
            .I(N__19652));
    Span4Mux_v I__1798 (
            .O(N__19652),
            .I(N__19649));
    Odrv4 I__1797 (
            .O(N__19649),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1796 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__1795 (
            .O(N__19643),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1794 (
            .O(N__19640),
            .I(N__19637));
    LocalMux I__1793 (
            .O(N__19637),
            .I(N__19634));
    Span4Mux_v I__1792 (
            .O(N__19634),
            .I(N__19631));
    Odrv4 I__1791 (
            .O(N__19631),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1790 (
            .O(N__19628),
            .I(N__19625));
    LocalMux I__1789 (
            .O(N__19625),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1788 (
            .O(N__19622),
            .I(N__19619));
    LocalMux I__1787 (
            .O(N__19619),
            .I(N__19616));
    Span4Mux_h I__1786 (
            .O(N__19616),
            .I(N__19613));
    Span4Mux_v I__1785 (
            .O(N__19613),
            .I(N__19610));
    Odrv4 I__1784 (
            .O(N__19610),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1783 (
            .O(N__19607),
            .I(N__19604));
    LocalMux I__1782 (
            .O(N__19604),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__1781 (
            .O(N__19601),
            .I(N__19598));
    LocalMux I__1780 (
            .O(N__19598),
            .I(N__19595));
    Span4Mux_v I__1779 (
            .O(N__19595),
            .I(N__19592));
    Odrv4 I__1778 (
            .O(N__19592),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1777 (
            .O(N__19589),
            .I(N__19586));
    LocalMux I__1776 (
            .O(N__19586),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__1775 (
            .O(N__19583),
            .I(N__19580));
    LocalMux I__1774 (
            .O(N__19580),
            .I(N__19577));
    Span4Mux_v I__1773 (
            .O(N__19577),
            .I(N__19574));
    Span4Mux_v I__1772 (
            .O(N__19574),
            .I(N__19571));
    Odrv4 I__1771 (
            .O(N__19571),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1770 (
            .O(N__19568),
            .I(N__19565));
    LocalMux I__1769 (
            .O(N__19565),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    CascadeMux I__1768 (
            .O(N__19562),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ));
    InMux I__1767 (
            .O(N__19559),
            .I(N__19553));
    InMux I__1766 (
            .O(N__19558),
            .I(N__19553));
    LocalMux I__1765 (
            .O(N__19553),
            .I(N__19550));
    Span4Mux_v I__1764 (
            .O(N__19550),
            .I(N__19547));
    Odrv4 I__1763 (
            .O(N__19547),
            .I(\pwm_generator_inst.O_10 ));
    CascadeMux I__1762 (
            .O(N__19544),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ));
    InMux I__1761 (
            .O(N__19541),
            .I(N__19538));
    LocalMux I__1760 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_v I__1759 (
            .O(N__19535),
            .I(N__19532));
    Span4Mux_v I__1758 (
            .O(N__19532),
            .I(N__19529));
    Odrv4 I__1757 (
            .O(N__19529),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1756 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__1755 (
            .O(N__19523),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1754 (
            .O(N__19520),
            .I(N__19517));
    LocalMux I__1753 (
            .O(N__19517),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__1752 (
            .O(N__19514),
            .I(N__19511));
    InMux I__1751 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__1750 (
            .O(N__19508),
            .I(N__19505));
    Span4Mux_v I__1749 (
            .O(N__19505),
            .I(N__19502));
    Span4Mux_v I__1748 (
            .O(N__19502),
            .I(N__19499));
    Odrv4 I__1747 (
            .O(N__19499),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1746 (
            .O(N__19496),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    CascadeMux I__1745 (
            .O(N__19493),
            .I(N__19490));
    InMux I__1744 (
            .O(N__19490),
            .I(N__19487));
    LocalMux I__1743 (
            .O(N__19487),
            .I(N__19484));
    Span4Mux_v I__1742 (
            .O(N__19484),
            .I(N__19481));
    Span4Mux_v I__1741 (
            .O(N__19481),
            .I(N__19478));
    Odrv4 I__1740 (
            .O(N__19478),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1739 (
            .O(N__19475),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1738 (
            .O(N__19472),
            .I(N__19469));
    LocalMux I__1737 (
            .O(N__19469),
            .I(N__19466));
    Span4Mux_v I__1736 (
            .O(N__19466),
            .I(N__19463));
    Span4Mux_v I__1735 (
            .O(N__19463),
            .I(N__19460));
    Odrv4 I__1734 (
            .O(N__19460),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1733 (
            .O(N__19457),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1732 (
            .O(N__19454),
            .I(N__19451));
    InMux I__1731 (
            .O(N__19451),
            .I(N__19448));
    LocalMux I__1730 (
            .O(N__19448),
            .I(N__19445));
    Span4Mux_v I__1729 (
            .O(N__19445),
            .I(N__19442));
    Span4Mux_v I__1728 (
            .O(N__19442),
            .I(N__19439));
    Odrv4 I__1727 (
            .O(N__19439),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1726 (
            .O(N__19436),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1725 (
            .O(N__19433),
            .I(N__19430));
    LocalMux I__1724 (
            .O(N__19430),
            .I(N__19427));
    Span4Mux_v I__1723 (
            .O(N__19427),
            .I(N__19424));
    Span4Mux_v I__1722 (
            .O(N__19424),
            .I(N__19421));
    Odrv4 I__1721 (
            .O(N__19421),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1720 (
            .O(N__19418),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1719 (
            .O(N__19415),
            .I(N__19412));
    InMux I__1718 (
            .O(N__19412),
            .I(N__19409));
    LocalMux I__1717 (
            .O(N__19409),
            .I(N__19406));
    Span4Mux_v I__1716 (
            .O(N__19406),
            .I(N__19403));
    Span4Mux_v I__1715 (
            .O(N__19403),
            .I(N__19400));
    Odrv4 I__1714 (
            .O(N__19400),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1713 (
            .O(N__19397),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1712 (
            .O(N__19394),
            .I(N__19391));
    LocalMux I__1711 (
            .O(N__19391),
            .I(N__19388));
    Span4Mux_v I__1710 (
            .O(N__19388),
            .I(N__19385));
    Span4Mux_v I__1709 (
            .O(N__19385),
            .I(N__19382));
    Odrv4 I__1708 (
            .O(N__19382),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1707 (
            .O(N__19379),
            .I(N__19375));
    InMux I__1706 (
            .O(N__19378),
            .I(N__19372));
    LocalMux I__1705 (
            .O(N__19375),
            .I(N__19369));
    LocalMux I__1704 (
            .O(N__19372),
            .I(N__19366));
    Span4Mux_v I__1703 (
            .O(N__19369),
            .I(N__19360));
    Span4Mux_h I__1702 (
            .O(N__19366),
            .I(N__19357));
    CascadeMux I__1701 (
            .O(N__19365),
            .I(N__19354));
    CascadeMux I__1700 (
            .O(N__19364),
            .I(N__19350));
    CascadeMux I__1699 (
            .O(N__19363),
            .I(N__19346));
    Span4Mux_v I__1698 (
            .O(N__19360),
            .I(N__19342));
    Span4Mux_v I__1697 (
            .O(N__19357),
            .I(N__19339));
    InMux I__1696 (
            .O(N__19354),
            .I(N__19326));
    InMux I__1695 (
            .O(N__19353),
            .I(N__19326));
    InMux I__1694 (
            .O(N__19350),
            .I(N__19326));
    InMux I__1693 (
            .O(N__19349),
            .I(N__19326));
    InMux I__1692 (
            .O(N__19346),
            .I(N__19326));
    InMux I__1691 (
            .O(N__19345),
            .I(N__19326));
    Odrv4 I__1690 (
            .O(N__19342),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    Odrv4 I__1689 (
            .O(N__19339),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    LocalMux I__1688 (
            .O(N__19326),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1687 (
            .O(N__19319),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1686 (
            .O(N__19316),
            .I(N__19313));
    LocalMux I__1685 (
            .O(N__19313),
            .I(N__19310));
    Odrv12 I__1684 (
            .O(N__19310),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1683 (
            .O(N__19307),
            .I(bfn_1_15_0_));
    InMux I__1682 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__1681 (
            .O(N__19301),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1680 (
            .O(N__19298),
            .I(N__19295));
    InMux I__1679 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__1678 (
            .O(N__19292),
            .I(N__19289));
    Span4Mux_v I__1677 (
            .O(N__19289),
            .I(N__19286));
    Span4Mux_v I__1676 (
            .O(N__19286),
            .I(N__19283));
    Odrv4 I__1675 (
            .O(N__19283),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    InMux I__1674 (
            .O(N__19280),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1673 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__1672 (
            .O(N__19274),
            .I(N__19271));
    Span4Mux_v I__1671 (
            .O(N__19271),
            .I(N__19268));
    Span4Mux_v I__1670 (
            .O(N__19268),
            .I(N__19265));
    Odrv4 I__1669 (
            .O(N__19265),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    CascadeMux I__1668 (
            .O(N__19262),
            .I(N__19259));
    InMux I__1667 (
            .O(N__19259),
            .I(N__19256));
    LocalMux I__1666 (
            .O(N__19256),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    InMux I__1665 (
            .O(N__19253),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1664 (
            .O(N__19250),
            .I(N__19247));
    LocalMux I__1663 (
            .O(N__19247),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1662 (
            .O(N__19244),
            .I(N__19241));
    InMux I__1661 (
            .O(N__19241),
            .I(N__19238));
    LocalMux I__1660 (
            .O(N__19238),
            .I(N__19235));
    Span4Mux_v I__1659 (
            .O(N__19235),
            .I(N__19232));
    Span4Mux_v I__1658 (
            .O(N__19232),
            .I(N__19229));
    Odrv4 I__1657 (
            .O(N__19229),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    InMux I__1656 (
            .O(N__19226),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1655 (
            .O(N__19223),
            .I(N__19220));
    LocalMux I__1654 (
            .O(N__19220),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1653 (
            .O(N__19217),
            .I(N__19214));
    InMux I__1652 (
            .O(N__19214),
            .I(N__19211));
    LocalMux I__1651 (
            .O(N__19211),
            .I(N__19208));
    Span4Mux_v I__1650 (
            .O(N__19208),
            .I(N__19205));
    Span4Mux_v I__1649 (
            .O(N__19205),
            .I(N__19202));
    Odrv4 I__1648 (
            .O(N__19202),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1647 (
            .O(N__19199),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1646 (
            .O(N__19196),
            .I(N__19193));
    LocalMux I__1645 (
            .O(N__19193),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__1644 (
            .O(N__19190),
            .I(N__19187));
    InMux I__1643 (
            .O(N__19187),
            .I(N__19184));
    LocalMux I__1642 (
            .O(N__19184),
            .I(N__19181));
    Span4Mux_v I__1641 (
            .O(N__19181),
            .I(N__19178));
    Span4Mux_v I__1640 (
            .O(N__19178),
            .I(N__19175));
    Odrv4 I__1639 (
            .O(N__19175),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    InMux I__1638 (
            .O(N__19172),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1637 (
            .O(N__19169),
            .I(N__19166));
    LocalMux I__1636 (
            .O(N__19166),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__1635 (
            .O(N__19163),
            .I(N__19160));
    InMux I__1634 (
            .O(N__19160),
            .I(N__19157));
    LocalMux I__1633 (
            .O(N__19157),
            .I(N__19154));
    Span4Mux_v I__1632 (
            .O(N__19154),
            .I(N__19151));
    Span4Mux_v I__1631 (
            .O(N__19151),
            .I(N__19148));
    Odrv4 I__1630 (
            .O(N__19148),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__1629 (
            .O(N__19145),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1628 (
            .O(N__19142),
            .I(N__19139));
    LocalMux I__1627 (
            .O(N__19139),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__1626 (
            .O(N__19136),
            .I(N__19133));
    InMux I__1625 (
            .O(N__19133),
            .I(N__19130));
    LocalMux I__1624 (
            .O(N__19130),
            .I(N__19127));
    Span4Mux_v I__1623 (
            .O(N__19127),
            .I(N__19124));
    Span4Mux_v I__1622 (
            .O(N__19124),
            .I(N__19121));
    Odrv4 I__1621 (
            .O(N__19121),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    InMux I__1620 (
            .O(N__19118),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1619 (
            .O(N__19115),
            .I(N__19112));
    LocalMux I__1618 (
            .O(N__19112),
            .I(N__19109));
    Odrv4 I__1617 (
            .O(N__19109),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__1616 (
            .O(N__19106),
            .I(N__19103));
    InMux I__1615 (
            .O(N__19103),
            .I(N__19100));
    LocalMux I__1614 (
            .O(N__19100),
            .I(N__19097));
    Span4Mux_v I__1613 (
            .O(N__19097),
            .I(N__19094));
    Span4Mux_v I__1612 (
            .O(N__19094),
            .I(N__19091));
    Odrv4 I__1611 (
            .O(N__19091),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    InMux I__1610 (
            .O(N__19088),
            .I(bfn_1_14_0_));
    InMux I__1609 (
            .O(N__19085),
            .I(N__19082));
    LocalMux I__1608 (
            .O(N__19082),
            .I(N__19079));
    Span4Mux_v I__1607 (
            .O(N__19079),
            .I(N__19076));
    Span4Mux_v I__1606 (
            .O(N__19076),
            .I(N__19073));
    Odrv4 I__1605 (
            .O(N__19073),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1604 (
            .O(N__19070),
            .I(N__19067));
    InMux I__1603 (
            .O(N__19067),
            .I(N__19064));
    LocalMux I__1602 (
            .O(N__19064),
            .I(N__19061));
    Odrv4 I__1601 (
            .O(N__19061),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1600 (
            .O(N__19058),
            .I(N__19054));
    InMux I__1599 (
            .O(N__19057),
            .I(N__19051));
    LocalMux I__1598 (
            .O(N__19054),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1597 (
            .O(N__19051),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    CascadeMux I__1596 (
            .O(N__19046),
            .I(N__19043));
    InMux I__1595 (
            .O(N__19043),
            .I(N__19040));
    LocalMux I__1594 (
            .O(N__19040),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_15_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_2_0_));
    defparam IN_MUX_bfv_15_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_3_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_15_3_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_15_28_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_12_11_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__23435),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_302_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNIEOIK_0  (
            .USERSIGNALTOGLOBALBUFFER(N__34529),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_181_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__29075),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_304_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__45908),
            .CLKHFEN(N__45912),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__45967),
            .RGB2PWM(N__19916),
            .RGB1(rgb_g),
            .CURREN(N__46081),
            .RGB2(rgb_b),
            .RGB1PWM(N__19910),
            .RGB0PWM(N__47925),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_6  (
            .in0(N__19379),
            .in1(N__21177),
            .in2(_gnd_net_),
            .in3(N__19057),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22700),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48482),
            .ce(),
            .sr(N__47816));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_6_3 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_6_3  (
            .in0(N__19058),
            .in1(N__19378),
            .in2(N__19046),
            .in3(N__21178),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2  (
            .in0(N__22400),
            .in1(N__21877),
            .in2(N__22699),
            .in3(N__22043),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48480),
            .ce(),
            .sr(N__47841));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_0 .LUT_INIT=16'b1000111110001100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_0  (
            .in0(N__22036),
            .in1(N__22136),
            .in2(N__22689),
            .in3(N__21873),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48476),
            .ce(),
            .sr(N__47850));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_1 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_1  (
            .in0(N__19946),
            .in1(N__20012),
            .in2(N__22217),
            .in3(N__22035),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48476),
            .ce(),
            .sr(N__47850));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_3  (
            .in0(N__20023),
            .in1(N__21974),
            .in2(N__20083),
            .in3(N__19960),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48476),
            .ce(),
            .sr(N__47850));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_4  (
            .in0(N__19959),
            .in1(N__20075),
            .in2(N__21053),
            .in3(N__20022),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48476),
            .ce(),
            .sr(N__47850));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_10_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_10_5  (
            .in0(N__20024),
            .in1(N__21983),
            .in2(N__20084),
            .in3(N__19961),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48476),
            .ce(),
            .sr(N__47850));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7 .LUT_INIT=16'b1101110011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7  (
            .in0(N__20082),
            .in1(N__20062),
            .in2(N__21878),
            .in3(N__20042),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48476),
            .ce(),
            .sr(N__47850));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_11_1 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_11_1  (
            .in0(N__22430),
            .in1(N__21870),
            .in2(N__22692),
            .in3(N__22039),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__47856));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_11_3 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_11_3  (
            .in0(N__22157),
            .in1(N__21869),
            .in2(N__22691),
            .in3(N__22038),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__47856));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7  (
            .in0(N__22181),
            .in1(N__21868),
            .in2(N__22690),
            .in3(N__22037),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__47856));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_12_2  (
            .in0(N__20296),
            .in1(N__21037),
            .in2(N__20324),
            .in3(N__21010),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_12_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__20134),
            .in2(_gnd_net_),
            .in3(N__19821),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__19085),
            .in2(N__19070),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__19304),
            .in2(N__19298),
            .in3(N__19280),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__19277),
            .in2(N__19262),
            .in3(N__19253),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__19250),
            .in2(N__19244),
            .in3(N__19226),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__19223),
            .in2(N__19217),
            .in3(N__19199),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__19196),
            .in2(N__19190),
            .in3(N__19172),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__19169),
            .in2(N__19163),
            .in3(N__19145),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__19142),
            .in2(N__19136),
            .in3(N__19118),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__19115),
            .in2(N__19106),
            .in3(N__19088),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__19520),
            .in2(N__19514),
            .in3(N__19496),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__19345),
            .in2(N__19493),
            .in3(N__19475),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__19472),
            .in2(N__19363),
            .in3(N__19457),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__19349),
            .in2(N__19454),
            .in3(N__19436),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__19433),
            .in2(N__19364),
            .in3(N__19418),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__19353),
            .in2(N__19415),
            .in3(N__19397),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__19394),
            .in2(N__19365),
            .in3(N__19319),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_15_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__19316),
            .in2(N__20417),
            .in3(N__19307),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_15_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_15_1 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_15_1  (
            .in0(N__19841),
            .in1(N__20693),
            .in2(N__19562),
            .in3(N__20675),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_15_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_15_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__20104),
            .in2(_gnd_net_),
            .in3(N__19786),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_1_15_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_1_15_7 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_1_15_7  (
            .in0(N__20141),
            .in1(N__19825),
            .in2(N__19802),
            .in3(N__20601),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_1_16_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_1_16_0 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_1_16_0  (
            .in0(N__20768),
            .in1(N__20749),
            .in2(N__19751),
            .in3(N__20598),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_16_1  (
            .in0(N__19873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19558),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_16_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_16_2  (
            .in0(N__19559),
            .in1(N__19859),
            .in2(N__19544),
            .in3(N__20596),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_16_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_16_4  (
            .in0(N__20732),
            .in1(N__20712),
            .in2(N__19736),
            .in3(N__20599),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_16_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_16_6  (
            .in0(N__20855),
            .in1(N__19934),
            .in2(N__20879),
            .in3(N__20600),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_1_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_1_16_7 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_1_16_7  (
            .in0(N__20597),
            .in1(N__20108),
            .in2(N__19766),
            .in3(N__19785),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__19526),
            .in2(_gnd_net_),
            .in3(N__19541),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__19706),
            .in2(_gnd_net_),
            .in3(N__19721),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__19688),
            .in2(_gnd_net_),
            .in3(N__19700),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__19667),
            .in2(_gnd_net_),
            .in3(N__19682),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__19646),
            .in2(_gnd_net_),
            .in3(N__19661),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__19628),
            .in2(_gnd_net_),
            .in3(N__19640),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__19607),
            .in2(_gnd_net_),
            .in3(N__19622),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__19589),
            .in2(_gnd_net_),
            .in3(N__19601),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__19568),
            .in2(_gnd_net_),
            .in3(N__19583),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__19883),
            .in2(_gnd_net_),
            .in3(N__19898),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__19877),
            .in2(_gnd_net_),
            .in3(N__19847),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_18_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_18_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_18_3  (
            .in0(N__20612),
            .in1(N__20192),
            .in2(_gnd_net_),
            .in3(N__19844),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_18_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__20667),
            .in2(_gnd_net_),
            .in3(N__19829),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_18_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__19826),
            .in2(_gnd_net_),
            .in3(N__19790),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_18_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__19787),
            .in2(_gnd_net_),
            .in3(N__19754),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_18_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__20748),
            .in2(_gnd_net_),
            .in3(N__19739),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__20714),
            .in2(_gnd_net_),
            .in3(N__19724),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_19_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20854),
            .in3(N__19925),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_19_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__20650),
            .in2(_gnd_net_),
            .in3(N__19922),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_19_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19919),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_1_29_3.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_29_3.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_29_3.LUT_INIT=16'b1100110000110011;
    LogicCell40 rgb_drv_RNO_0_LC_1_29_3 (
            .in0(_gnd_net_),
            .in1(N__45541),
            .in2(_gnd_net_),
            .in3(N__47923),
            .lcout(N_34_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_1_30_0.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_1_30_0.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_1_30_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_1_30_0 (
            .in0(N__47924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45545),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_8_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_2_9_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19904),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48477),
            .ce(),
            .sr(N__47832));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24746),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48477),
            .ce(),
            .sr(N__47832));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_2_9_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_2_9_7 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_2_9_7  (
            .in0(N__21323),
            .in1(N__21408),
            .in2(N__21269),
            .in3(N__20810),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48477),
            .ce(),
            .sr(N__47832));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_10_0 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_10_0  (
            .in0(N__22209),
            .in1(N__22667),
            .in2(_gnd_net_),
            .in3(N__20337),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__22208),
            .in2(_gnd_net_),
            .in3(N__20058),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_10_4 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_10_4  (
            .in0(N__22669),
            .in1(N__19945),
            .in2(N__20087),
            .in3(N__22034),
            .lcout(\current_shift_inst.PI_CTRL.N_166 ),
            .ltout(\current_shift_inst.PI_CTRL.N_166_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_10_5 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_10_5  (
            .in0(N__20063),
            .in1(N__20038),
            .in2(N__20027),
            .in3(N__21871),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6  (
            .in0(N__21872),
            .in1(N__22668),
            .in2(N__22216),
            .in3(N__20338),
            .lcout(\current_shift_inst.PI_CTRL.N_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_7  (
            .in0(N__20005),
            .in1(N__19990),
            .in2(_gnd_net_),
            .in3(N__19975),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_11_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_11_0  (
            .in0(N__22673),
            .in1(N__20339),
            .in2(_gnd_net_),
            .in3(N__21867),
            .lcout(\current_shift_inst.PI_CTRL.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_11_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_11_1  (
            .in0(N__22429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22176),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_11_2  (
            .in0(N__22132),
            .in1(N__22393),
            .in2(N__19949),
            .in3(N__22156),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_2_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_2_11_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__22428),
            .in2(_gnd_net_),
            .in3(N__22155),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_7  (
            .in0(N__22392),
            .in1(N__22131),
            .in2(N__20342),
            .in3(N__22177),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_12_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_12_2  (
            .in0(N__20266),
            .in1(N__20323),
            .in2(N__20990),
            .in3(N__20297),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_12_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_12_3 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_12_3  (
            .in0(N__20279),
            .in1(N__20247),
            .in2(N__20270),
            .in3(N__20215),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_12_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_12_5  (
            .in0(N__20267),
            .in1(N__20248),
            .in2(N__20225),
            .in3(N__20216),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__20191),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__20168),
            .in2(_gnd_net_),
            .in3(N__20156),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__20153),
            .in2(_gnd_net_),
            .in3(N__20123),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__20120),
            .in2(_gnd_net_),
            .in3(N__20090),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__20408),
            .in2(_gnd_net_),
            .in3(N__20402),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__45836),
            .in2(N__20399),
            .in3(N__20390),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__20387),
            .in2(N__45889),
            .in3(N__20381),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__20378),
            .in2(N__45856),
            .in3(N__20372),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__20369),
            .in2(_gnd_net_),
            .in3(N__20363),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__20360),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__20354),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__20348),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__20468),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__20462),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__20456),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__20450),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__20444),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__20438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__20432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__20426),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_15_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20420),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__20543),
            .in2(N__20617),
            .in3(N__20611),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__20537),
            .in2(_gnd_net_),
            .in3(N__20528),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__20525),
            .in2(_gnd_net_),
            .in3(N__20519),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_16_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20516),
            .in3(N__20507),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__20504),
            .in2(_gnd_net_),
            .in3(N__20498),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__20495),
            .in2(_gnd_net_),
            .in3(N__20489),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__20486),
            .in2(_gnd_net_),
            .in3(N__20480),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__20477),
            .in2(_gnd_net_),
            .in3(N__20471),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_17_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20552),
            .in3(N__20795),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_17_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_17_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_17_1  (
            .in0(N__20792),
            .in1(N__20616),
            .in2(N__20783),
            .in3(N__20771),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_4  (
            .in0(N__20750),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20767),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_5  (
            .in0(N__20713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20731),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_17_6  (
            .in0(N__20671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20692),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_18_1  (
            .in0(N__20651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20638),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_18_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_18_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_18_2  (
            .in0(N__20639),
            .in1(N__20627),
            .in2(N__20621),
            .in3(N__20618),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_2_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_2_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_2_18_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_2_18_5  (
            .in0(N__34008),
            .in1(N__34284),
            .in2(N__33592),
            .in3(N__34183),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48405),
            .ce(N__28847),
            .sr(N__47882));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_2_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_2_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_2_18_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_2_18_6  (
            .in0(N__34184),
            .in1(N__33703),
            .in2(N__34336),
            .in3(N__34009),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48405),
            .ce(N__28847),
            .sr(N__47882));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_19_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_19_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__20872),
            .in2(_gnd_net_),
            .in3(N__20853),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_21_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_21_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_21_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_3_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_3_8_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNITBL3_9_LC_3_8_0  (
            .in0(N__21923),
            .in1(N__21530),
            .in2(_gnd_net_),
            .in3(N__21640),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_3_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_3_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIRPD2_0_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(N__21093),
            .in2(_gnd_net_),
            .in3(N__21069),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_3_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_3_8_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_2_LC_3_8_4  (
            .in0(N__21673),
            .in1(N__21712),
            .in2(N__20831),
            .in3(N__21748),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_3_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_3_8_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_6_LC_3_8_5  (
            .in0(N__20828),
            .in1(N__21568),
            .in2(N__20822),
            .in3(N__21617),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_3_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_3_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_3_9_0  (
            .in0(N__20927),
            .in1(N__21095),
            .in2(_gnd_net_),
            .in3(N__20819),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_1_LC_3_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_3_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_3_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_3_9_1  (
            .in0(N__20912),
            .in1(N__21071),
            .in2(_gnd_net_),
            .in3(N__20816),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_2_LC_3_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_3_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_3_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_3_9_2  (
            .in0(N__20928),
            .in1(N__21749),
            .in2(_gnd_net_),
            .in3(N__20813),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_3_LC_3_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_3_9_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_3_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_3_9_3  (
            .in0(N__20913),
            .in1(N__21713),
            .in2(_gnd_net_),
            .in3(N__20948),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_4_LC_3_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_3_9_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_3_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_3_9_4  (
            .in0(N__20929),
            .in1(N__21674),
            .in2(_gnd_net_),
            .in3(N__20945),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_5_LC_3_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_3_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_3_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_3_9_5  (
            .in0(N__20914),
            .in1(N__21641),
            .in2(_gnd_net_),
            .in3(N__20942),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_6_LC_3_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_3_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_3_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_3_9_6  (
            .in0(N__20930),
            .in1(N__21616),
            .in2(_gnd_net_),
            .in3(N__20939),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_7_LC_3_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_3_9_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_3_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_3_9_7  (
            .in0(N__20915),
            .in1(N__21569),
            .in2(_gnd_net_),
            .in3(N__20936),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__48475),
            .ce(),
            .sr(N__47823));
    defparam \pwm_generator_inst.counter_8_LC_3_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_3_10_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_3_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_3_10_0  (
            .in0(N__20926),
            .in1(N__21529),
            .in2(_gnd_net_),
            .in3(N__20933),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__48469),
            .ce(),
            .sr(N__47833));
    defparam \pwm_generator_inst.counter_9_LC_3_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_3_10_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_3_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_9_LC_3_10_1  (
            .in0(N__20925),
            .in1(N__21922),
            .in2(_gnd_net_),
            .in3(N__20882),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(),
            .sr(N__47833));
    defparam \pwm_generator_inst.threshold_6_LC_3_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_3_10_2 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_3_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21482),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(),
            .sr(N__47833));
    defparam \pwm_generator_inst.threshold_5_LC_3_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_3_10_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_3_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21443),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(),
            .sr(N__47833));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23750),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48462),
            .ce(),
            .sr(N__47842));
    defparam \pwm_generator_inst.threshold_3_LC_3_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_3_11_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_3_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21497),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48462),
            .ce(),
            .sr(N__47842));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_12_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(N__21038),
            .in2(_gnd_net_),
            .in3(N__21014),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_0_LC_3_13_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_3_13_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_3_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20957),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48443),
            .ce(),
            .sr(N__47857));
    defparam \pwm_generator_inst.threshold_7_LC_3_13_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_3_13_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_3_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20972),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48443),
            .ce(),
            .sr(N__47857));
    defparam \pwm_generator_inst.threshold_9_LC_3_14_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_3_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21428),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48434),
            .ce(),
            .sr(N__47862));
    defparam \pwm_generator_inst.threshold_4_LC_3_14_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_3_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21464),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48434),
            .ce(),
            .sr(N__47862));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_15_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_15_2 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_15_2 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_15_2  (
            .in0(N__21253),
            .in1(N__21407),
            .in2(N__21348),
            .in3(N__20978),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48425),
            .ce(),
            .sr(N__47869));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_15_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_15_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_3_15_5  (
            .in0(N__21404),
            .in1(N__20963),
            .in2(N__21346),
            .in3(N__21254),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48425),
            .ce(),
            .sr(N__47869));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_15_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_15_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_15_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_3_15_6  (
            .in0(N__21252),
            .in1(N__21406),
            .in2(N__21347),
            .in3(N__21503),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48425),
            .ce(),
            .sr(N__47869));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_15_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_15_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_15_7 .LUT_INIT=16'b1111111100110101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_3_15_7  (
            .in0(N__21405),
            .in1(N__21330),
            .in2(N__21273),
            .in3(N__21488),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48425),
            .ce(),
            .sr(N__47869));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_16_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_3_16_2  (
            .in0(N__21410),
            .in1(N__21289),
            .in2(N__21359),
            .in3(N__21470),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48413),
            .ce(),
            .sr(N__47873));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_16_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_16_4 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_3_16_4  (
            .in0(N__21409),
            .in1(N__21455),
            .in2(N__21358),
            .in3(N__21288),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48413),
            .ce(),
            .sr(N__47873));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_16_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_16_5 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_3_16_5  (
            .in0(N__21286),
            .in1(N__21355),
            .in2(N__21418),
            .in3(N__21449),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48413),
            .ce(),
            .sr(N__47873));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_16_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_16_7 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_3_16_7  (
            .in0(N__21287),
            .in1(N__21356),
            .in2(N__21419),
            .in3(N__21434),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48413),
            .ce(),
            .sr(N__47873));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_17_6 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_3_17_6  (
            .in0(N__21411),
            .in1(N__21357),
            .in2(N__21290),
            .in3(N__21116),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48406),
            .ce(),
            .sr(N__47877));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__21077),
            .in2(N__21110),
            .in3(N__21094),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__21755),
            .in2(N__21800),
            .in3(N__21070),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_9_2  (
            .in0(N__21747),
            .in1(N__21731),
            .in2(N__21779),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__21695),
            .in2(N__21725),
            .in3(N__21711),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__21656),
            .in2(N__21689),
            .in3(N__21672),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__21623),
            .in2(N__21650),
            .in3(N__21639),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_9_6  (
            .in0(N__21615),
            .in1(N__21590),
            .in2(N__21599),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__21551),
            .in2(N__21584),
            .in3(N__21567),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__21509),
            .in2(N__21545),
            .in3(N__21528),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__21902),
            .in2(N__21938),
            .in3(N__21921),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_4_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_4_10_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_4_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21896),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48463),
            .ce(),
            .sr(N__47824));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_13_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_13_1  (
            .in0(N__21962),
            .in1(N__21812),
            .in2(N__21956),
            .in3(N__22073),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_4_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_4_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__22741),
            .in2(_gnd_net_),
            .in3(N__22363),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_4_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_4_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_4_14_3  (
            .in0(N__22721),
            .in1(N__22766),
            .in2(N__21815),
            .in3(N__22787),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_1_LC_4_15_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_4_15_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_4_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21806),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48414),
            .ce(),
            .sr(N__47863));
    defparam \pwm_generator_inst.threshold_2_LC_4_15_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_4_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21788),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48414),
            .ce(),
            .sr(N__47863));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_8_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_8_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21764),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48470),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_5_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_5_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27567),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24782),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(),
            .sr(N__47817));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23516),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(),
            .sr(N__47817));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_5_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_5_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27723),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_5_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_5_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28464),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_5_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_5_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_5_12_0  (
            .in0(N__22240),
            .in1(N__22255),
            .in2(N__22597),
            .in3(N__22270),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_5_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_5_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_5_12_3  (
            .in0(N__22559),
            .in1(N__22574),
            .in2(N__22601),
            .in3(N__22241),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_5_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_5_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_5_12_4  (
            .in0(N__22294),
            .in1(N__22256),
            .in2(N__22336),
            .in3(N__22271),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_5_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_5_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_5_12_5  (
            .in0(N__22537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22519),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_5_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_5_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_5_12_6  (
            .in0(N__22573),
            .in1(N__22558),
            .in2(N__21947),
            .in3(N__21944),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_5_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_5_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_5_13_0  (
            .in0(N__22295),
            .in1(N__22745),
            .in2(N__22460),
            .in3(N__22364),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_5_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_5_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__22831),
            .in2(_gnd_net_),
            .in3(N__22495),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_5_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_5_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_5_13_2  (
            .in0(N__22477),
            .in1(N__22802),
            .in2(N__22085),
            .in3(N__22817),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_5_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_5_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__22801),
            .in2(_gnd_net_),
            .in3(N__22816),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_5_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_5_13_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_5_13_6  (
            .in0(N__22496),
            .in1(N__22520),
            .in2(N__22481),
            .in3(N__22541),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_5_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_5_13_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_5_13_7  (
            .in0(N__22459),
            .in1(N__22832),
            .in2(N__22082),
            .in3(N__22079),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_5_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_5_14_2  (
            .in0(N__22762),
            .in1(N__22786),
            .in2(N__22337),
            .in3(N__22720),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_5_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_5_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_5_14_3  (
            .in0(N__22067),
            .in1(N__22061),
            .in2(N__22052),
            .in3(N__22049),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_14_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_14_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_5_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21995),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48415),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_5_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_5_20_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_5_20_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_5_20_4  (
            .in0(N__33524),
            .in1(N__23051),
            .in2(_gnd_net_),
            .in3(N__33141),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48380),
            .ce(),
            .sr(N__47879));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_2_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_2_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22109),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48481),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_4_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_4_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22100),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48478),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_7_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_7_8_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_7_8_6  (
            .in0(N__28298),
            .in1(N__28094),
            .in2(_gnd_net_),
            .in3(N__25196),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48453),
            .ce(),
            .sr(N__47798));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_7_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_7_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__31185),
            .in2(_gnd_net_),
            .in3(N__31601),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_9_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__23704),
            .in2(_gnd_net_),
            .in3(N__24935),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_9_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_9_2  (
            .in0(N__24965),
            .in1(N__24880),
            .in2(N__22091),
            .in3(N__27297),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_9_3 .LUT_INIT=16'b1111001011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_9_3  (
            .in0(N__23096),
            .in1(N__23656),
            .in2(N__22088),
            .in3(N__24745),
            .lcout(\current_shift_inst.PI_CTRL.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_7_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_7_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_7_9_5  (
            .in0(N__31600),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27406),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_7_10_1  (
            .in0(N__29696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48435),
            .ce(),
            .sr(N__47807));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29770),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48435),
            .ce(),
            .sr(N__47807));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29860),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48435),
            .ce(),
            .sr(N__47807));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27017),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48435),
            .ce(),
            .sr(N__47807));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__29818),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48435),
            .ce(),
            .sr(N__47807));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__23660),
            .in2(N__22226),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__24934),
            .in2(N__23606),
            .in3(N__22160),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__27302),
            .in2(N__23621),
            .in3(N__22139),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__23705),
            .in2(N__23765),
            .in3(N__22112),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__24976),
            .in2(N__22439),
            .in3(N__22412),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__24886),
            .in2(N__22409),
            .in3(N__22376),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__25024),
            .in2(N__22373),
            .in3(N__22340),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__31919),
            .in2(N__24797),
            .in3(N__22307),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__48426),
            .ce(),
            .sr(N__47812));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__22304),
            .in2(N__31616),
            .in3(N__22274),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__31267),
            .in2(N__29990),
            .in3(N__22259),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__31189),
            .in2(N__29948),
            .in3(N__22244),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__27402),
            .in2(N__23717),
            .in3(N__22229),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__28471),
            .in2(N__28633),
            .in3(N__22577),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__28602),
            .in2(N__27574),
            .in3(N__22562),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__31740),
            .in2(N__28634),
            .in3(N__22544),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__28606),
            .in2(N__31796),
            .in3(N__22523),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__48416),
            .ce(),
            .sr(N__47818));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__29516),
            .in2(N__28659),
            .in3(N__22499),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__28638),
            .in2(N__31855),
            .in3(N__22484),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__31685),
            .in2(N__28660),
            .in3(N__22463),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__28642),
            .in2(N__27461),
            .in3(N__22442),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__27724),
            .in2(N__28661),
            .in3(N__22820),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__28646),
            .in2(N__27645),
            .in3(N__22805),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__28725),
            .in2(N__28662),
            .in3(N__22790),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__28650),
            .in2(N__27226),
            .in3(N__22769),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__48407),
            .ce(),
            .sr(N__47825));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__28397),
            .in2(N__28663),
            .in3(N__22748),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__48399),
            .ce(),
            .sr(N__47834));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__28654),
            .in2(N__28352),
            .in3(N__22724),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__48399),
            .ce(),
            .sr(N__47834));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__27772),
            .in2(N__28664),
            .in3(N__22706),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__48399),
            .ce(),
            .sr(N__47834));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_14_3  (
            .in0(N__27903),
            .in1(N__28658),
            .in2(_gnd_net_),
            .in3(N__22703),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48399),
            .ce(),
            .sr(N__47834));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__22880),
            .in2(N__23162),
            .in3(N__23868),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__22874),
            .in2(N__23327),
            .in3(N__23851),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__22868),
            .in2(N__23150),
            .in3(N__23830),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__22862),
            .in2(N__23315),
            .in3(N__23806),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__22856),
            .in2(N__23303),
            .in3(N__23785),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__22850),
            .in2(N__23189),
            .in3(N__24061),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_15_7  (
            .in0(N__24040),
            .in1(N__22844),
            .in2(N__23288),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_16_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_16_0  (
            .in0(N__24020),
            .in1(N__22838),
            .in2(N__23273),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__22964),
            .in2(N__23177),
            .in3(N__23996),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_16_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_16_2  (
            .in0(N__23971),
            .in1(N__22940),
            .in2(N__22958),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__22916),
            .in2(N__22934),
            .in3(N__23950),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__22910),
            .in2(N__22991),
            .in3(N__23929),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__22904),
            .in2(N__23234),
            .in3(N__23908),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__22898),
            .in2(N__23264),
            .in3(N__24187),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__22892),
            .in2(N__23336),
            .in3(N__24166),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__22886),
            .in2(N__28859),
            .in3(N__25940),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__23036),
            .in2(N__23015),
            .in3(N__24143),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_17_2  (
            .in0(N__24119),
            .in1(N__23030),
            .in2(N__23003),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__23024),
            .in2(N__28874),
            .in3(N__24095),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23018),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__25979),
            .in2(_gnd_net_),
            .in3(N__35601),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_18_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_7_18_2  (
            .in0(N__30230),
            .in1(N__33992),
            .in2(_gnd_net_),
            .in3(N__34360),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48381),
            .ce(N__28842),
            .sr(N__47864));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_18_3 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__34357),
            .in2(N__34010),
            .in3(N__30770),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48381),
            .ce(N__28842),
            .sr(N__47864));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_7_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_7_18_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_7_18_5  (
            .in0(N__34359),
            .in1(N__33743),
            .in2(N__34012),
            .in3(N__34177),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48381),
            .ce(N__28842),
            .sr(N__47864));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_7  (
            .in0(N__34358),
            .in1(N__34176),
            .in2(N__34011),
            .in3(N__32569),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48381),
            .ce(N__28842),
            .sr(N__47864));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_7_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_7_19_3 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_7_19_3  (
            .in0(N__33514),
            .in1(N__23366),
            .in2(_gnd_net_),
            .in3(N__33142),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48376),
            .ce(),
            .sr(N__47870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25922),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48371),
            .ce(N__24595),
            .sr(N__47874));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25889),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48371),
            .ce(N__24595),
            .sr(N__47874));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_7_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_7_21_0 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_7_21_0  (
            .in0(N__24391),
            .in1(N__24241),
            .in2(N__24521),
            .in3(N__29053),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_10_LC_7_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_10_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_10_LC_7_21_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_10_LC_7_21_1  (
            .in0(N__33585),
            .in1(N__24392),
            .in2(_gnd_net_),
            .in3(N__33203),
            .lcout(\delay_measurement_inst.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI53F91_1_LC_7_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI53F91_1_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI53F91_1_LC_7_21_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI53F91_1_LC_7_21_2  (
            .in0(N__24220),
            .in1(N__29052),
            .in2(_gnd_net_),
            .in3(N__26680),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_7_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_7_21_3 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_7_21_3  (
            .in0(N__24242),
            .in1(N__30487),
            .in2(N__23039),
            .in3(N__24484),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_19_LC_7_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_19_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_19_LC_7_21_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_19_LC_7_21_4  (
            .in0(N__33205),
            .in1(N__30285),
            .in2(_gnd_net_),
            .in3(N__24520),
            .lcout(\delay_measurement_inst.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_8_LC_7_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_8_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_8_LC_7_21_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_8_LC_7_21_5  (
            .in0(N__24428),
            .in1(N__32659),
            .in2(_gnd_net_),
            .in3(N__33206),
            .lcout(\delay_measurement_inst.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_11_LC_7_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_11_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_11_LC_7_21_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_11_LC_7_21_7  (
            .in0(N__33685),
            .in1(N__24368),
            .in2(_gnd_net_),
            .in3(N__33204),
            .lcout(\delay_measurement_inst.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_7_22_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_7_22_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_7_22_0  (
            .in0(N__33452),
            .in1(N__23081),
            .in2(_gnd_net_),
            .in3(N__33132),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48359),
            .ce(),
            .sr(N__47880));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_7_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_7_22_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_7_22_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_7_22_4  (
            .in0(N__33451),
            .in1(N__23075),
            .in2(_gnd_net_),
            .in3(N__33131),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48359),
            .ce(),
            .sr(N__47880));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_7_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_7_23_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_7_23_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_7_23_1  (
            .in0(N__33138),
            .in1(N__33509),
            .in2(_gnd_net_),
            .in3(N__23069),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48353),
            .ce(),
            .sr(N__47883));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_7_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_7_23_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_7_23_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_7_23_5  (
            .in0(N__33136),
            .in1(N__33507),
            .in2(_gnd_net_),
            .in3(N__23420),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48353),
            .ce(),
            .sr(N__47883));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_7_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_7_23_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_7_23_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_7_23_7  (
            .in0(N__33137),
            .in1(N__33508),
            .in2(_gnd_net_),
            .in3(N__23441),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48353),
            .ce(),
            .sr(N__47883));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_3_5 (
            .in0(N__23060),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48479),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_8_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_8_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_8_6_5 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst2.state_0_LC_8_6_5  (
            .in0(N__23541),
            .in1(N__38000),
            .in2(N__23575),
            .in3(N__23591),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48464),
            .ce(),
            .sr(N__47788));
    defparam \phase_controller_inst2.state_1_LC_8_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_8_7_5 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst2.state_1_LC_8_7_5  (
            .in0(N__35762),
            .in1(N__23543),
            .in2(N__23574),
            .in3(N__36818),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48454),
            .ce(),
            .sr(N__47791));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_8_0 .LUT_INIT=16'b0000000111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_8_8_0  (
            .in0(N__28301),
            .in1(N__27967),
            .in2(N__28132),
            .in3(N__25448),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(N__47795));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_8_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_8_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_8_8_3  (
            .in0(N__31739),
            .in1(N__25017),
            .in2(N__23222),
            .in3(N__23480),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_8_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_8_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_8_8_4  (
            .in0(N__23129),
            .in1(N__23105),
            .in2(N__23111),
            .in3(N__23138),
            .lcout(\current_shift_inst.PI_CTRL.N_74 ),
            .ltout(\current_shift_inst.PI_CTRL.N_74_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_8_5 .LUT_INIT=16'b0000000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_8_8_5  (
            .in0(N__27966),
            .in1(N__28302),
            .in2(N__23108),
            .in3(N__25409),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(N__47795));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36740),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36725),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36689),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_8_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_8_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29691),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_8_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_8_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30013),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_10_0  (
            .in0(N__31846),
            .in1(N__28396),
            .in2(N__27649),
            .in3(N__28729),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_1  (
            .in0(N__24778),
            .in1(N__23514),
            .in2(_gnd_net_),
            .in3(N__23743),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_8_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_8_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_8_10_2  (
            .in0(N__27219),
            .in1(N__27765),
            .in2(N__23090),
            .in3(N__23120),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_8_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_8_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24885),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_10_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__24969),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_8_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_8_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_8_10_6  (
            .in0(N__27707),
            .in1(N__31678),
            .in2(N__31785),
            .in3(N__27885),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27641),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_8_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_8_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23698),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_8_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_8_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_8_11_2  (
            .in0(N__27442),
            .in1(N__28450),
            .in2(N__28351),
            .in3(N__31250),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_8_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_8_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_8_11_3  (
            .in0(N__28347),
            .in1(N__27443),
            .in2(N__27914),
            .in3(N__25009),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_8_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_8_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31249),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_11_7  (
            .in0(N__27550),
            .in1(N__27391),
            .in2(N__29503),
            .in3(N__31918),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI764B_28_LC_8_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI764B_28_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI764B_28_LC_8_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI764B_28_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__28392),
            .in2(_gnd_net_),
            .in3(N__31611),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_29_LC_8_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_29_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_29_LC_8_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_29_LC_8_12_5  (
            .in0(N__23474),
            .in1(N__23210),
            .in2(N__30971),
            .in3(N__23204),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(\current_shift_inst.PI_CTRL.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_12_6 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_8_12_6  (
            .in0(N__27886),
            .in1(N__28144),
            .in2(N__23192),
            .in3(N__25703),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48408),
            .ce(),
            .sr(N__47813));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_8_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_8_13_0 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_8_13_0  (
            .in0(N__34155),
            .in1(N__34004),
            .in2(N__30452),
            .in3(N__34340),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(N__28831),
            .sr(N__47819));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_8_13_1 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_8_13_1  (
            .in0(N__34339),
            .in1(N__33643),
            .in2(N__34013),
            .in3(N__34156),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(N__28831),
            .sr(N__47819));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_8_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_8_13_5 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_8_13_5  (
            .in0(N__34002),
            .in1(N__32875),
            .in2(_gnd_net_),
            .in3(N__32818),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(N__28831),
            .sr(N__47819));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_8_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_8_13_6 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_8_13_6  (
            .in0(N__32819),
            .in1(N__34003),
            .in2(_gnd_net_),
            .in3(N__32795),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(N__28831),
            .sr(N__47819));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_14_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_14_0  (
            .in0(N__35543),
            .in1(N__35425),
            .in2(N__35325),
            .in3(N__24029),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48395),
            .ce(),
            .sr(N__47826));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_14_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_14_1  (
            .in0(N__35424),
            .in1(N__35545),
            .in2(N__35324),
            .in3(N__24005),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48395),
            .ce(),
            .sr(N__47826));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_2  (
            .in0(N__35544),
            .in1(N__35426),
            .in2(N__35326),
            .in3(N__23981),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48395),
            .ce(),
            .sr(N__47826));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_14_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_14_4  (
            .in0(N__35542),
            .in1(N__35291),
            .in2(_gnd_net_),
            .in3(N__35423),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0  (
            .in0(N__35308),
            .in1(N__35431),
            .in2(N__35578),
            .in3(N__24128),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1  (
            .in0(N__35427),
            .in1(N__35546),
            .in2(N__35327),
            .in3(N__24104),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2  (
            .in0(N__35309),
            .in1(N__35432),
            .in2(N__35579),
            .in3(N__24077),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_15_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_15_3  (
            .in0(N__35428),
            .in1(N__35547),
            .in2(N__35328),
            .in3(N__23840),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_15_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_15_4  (
            .in0(N__35310),
            .in1(N__35433),
            .in2(N__35580),
            .in3(N__23819),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_15_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_15_5  (
            .in0(N__35429),
            .in1(N__35548),
            .in2(N__35329),
            .in3(N__23795),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_15_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_15_6  (
            .in0(N__35311),
            .in1(N__35434),
            .in2(N__35581),
            .in3(N__23774),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_15_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_15_7  (
            .in0(N__35430),
            .in1(N__35549),
            .in2(N__35330),
            .in3(N__24050),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(N__47835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_16_0 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_16_0  (
            .in0(N__35301),
            .in1(N__23960),
            .in2(N__35584),
            .in3(N__35440),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_8_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_8_16_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_8_16_1  (
            .in0(N__25978),
            .in1(N__23872),
            .in2(_gnd_net_),
            .in3(N__35609),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_16_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_16_2  (
            .in0(N__35304),
            .in1(N__35527),
            .in2(N__23237),
            .in3(N__35441),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_16_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_16_3  (
            .in0(N__35435),
            .in1(N__35305),
            .in2(N__35571),
            .in3(N__23939),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_16_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_16_4  (
            .in0(N__35302),
            .in1(N__35438),
            .in2(N__35582),
            .in3(N__23918),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_16_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_16_5  (
            .in0(N__35436),
            .in1(N__35306),
            .in2(N__35572),
            .in3(N__23897),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_16_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_16_6  (
            .in0(N__35303),
            .in1(N__35439),
            .in2(N__35583),
            .in3(N__24176),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_16_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_16_7  (
            .in0(N__35437),
            .in1(N__35307),
            .in2(N__35573),
            .in3(N__24155),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(),
            .sr(N__47843));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_8_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_8_17_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_8_17_0  (
            .in0(N__33945),
            .in1(N__34341),
            .in2(N__34506),
            .in3(N__34097),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_8_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_8_17_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_8_17_1  (
            .in0(N__34099),
            .in1(N__34424),
            .in2(N__34362),
            .in3(N__33956),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_8_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_8_17_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_8_17_2  (
            .in0(N__33946),
            .in1(N__34100),
            .in2(N__34058),
            .in3(N__34356),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_8_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_8_17_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_8_17_3  (
            .in0(N__34101),
            .in1(N__33947),
            .in2(N__34363),
            .in3(N__32431),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_8_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_8_17_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_8_17_4  (
            .in0(N__32369),
            .in1(N__34342),
            .in2(N__33985),
            .in3(N__34102),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_8_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_8_17_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_8_17_5  (
            .in0(N__34103),
            .in1(N__33948),
            .in2(N__34364),
            .in3(N__32724),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_17_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_8_17_6  (
            .in0(N__32670),
            .in1(N__34343),
            .in2(N__33986),
            .in3(N__34104),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_17_7 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_8_17_7  (
            .in0(N__34098),
            .in1(N__30362),
            .in2(N__34361),
            .in3(N__33955),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48382),
            .ce(N__28832),
            .sr(N__47851));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_8_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_8_18_1 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_8_18_1  (
            .in0(N__33140),
            .in1(N__23372),
            .in2(N__33523),
            .in3(_gnd_net_),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48377),
            .ce(),
            .sr(N__47858));
    defparam \phase_controller_inst2.S2_LC_8_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.S2_LC_8_18_4  (
            .in0(N__23579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48377),
            .ce(),
            .sr(N__47858));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_8_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_8_18_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_8_18_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_8_18_6  (
            .in0(N__24254),
            .in1(N__33500),
            .in2(_gnd_net_),
            .in3(N__33139),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48377),
            .ce(),
            .sr(N__47858));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_7_LC_8_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_7_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_7_LC_8_19_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_7_LC_8_19_0  (
            .in0(N__33273),
            .in1(N__32723),
            .in2(_gnd_net_),
            .in3(N__24450),
            .lcout(\delay_measurement_inst.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_19_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_19_2  (
            .in0(N__24414),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24449),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_16_LC_8_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_16_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_16_LC_8_19_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_16_LC_8_19_6  (
            .in0(N__33272),
            .in1(_gnd_net_),
            .in2(N__32920),
            .in3(N__24571),
            .lcout(\delay_measurement_inst.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_14_LC_8_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_14_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_14_LC_8_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_14_LC_8_19_7  (
            .in0(N__30349),
            .in1(N__24287),
            .in2(_gnd_net_),
            .in3(N__33271),
            .lcout(\delay_measurement_inst.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_20_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_20_1  (
            .in0(N__24304),
            .in1(N__24361),
            .in2(N__24337),
            .in3(N__24385),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFRS4_9_LC_8_20_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFRS4_9_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFRS4_9_LC_8_20_2 .LUT_INIT=16'b0101000011010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFRS4_9_LC_8_20_2  (
            .in0(N__28758),
            .in1(N__23360),
            .in2(N__23354),
            .in3(N__23351),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_8_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_8_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_8_20_3  (
            .in0(N__24303),
            .in1(N__28757),
            .in2(N__24572),
            .in3(N__24471),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_20_4  (
            .in0(N__24546),
            .in1(N__24516),
            .in2(N__28977),
            .in3(N__24570),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JGD6_14_LC_8_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JGD6_14_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JGD6_14_LC_8_20_5 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JGD6_14_LC_8_20_5  (
            .in0(N__26764),
            .in1(N__24286),
            .in2(N__23345),
            .in3(N__23342),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_20_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_20_6  (
            .in0(N__24472),
            .in1(N__24415),
            .in2(_gnd_net_),
            .in3(N__24451),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_8_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_8_20_7 .LUT_INIT=16'b0100110001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_8_20_7  (
            .in0(N__23414),
            .in1(N__24285),
            .in2(N__23408),
            .in3(N__28759),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_4_LC_8_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_4_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_4_LC_8_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_4_LC_8_21_0  (
            .in0(N__24219),
            .in1(N__32426),
            .in2(_gnd_net_),
            .in3(N__33202),
            .lcout(\delay_measurement_inst.N_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_8_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_8_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_8_21_1  (
            .in0(N__24284),
            .in1(N__24360),
            .in2(N__24336),
            .in3(N__26762),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJAU73_7_LC_8_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJAU73_7_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJAU73_7_LC_8_21_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJAU73_7_LC_8_21_2  (
            .in0(N__24427),
            .in1(N__24455),
            .in2(N__23405),
            .in3(N__23402),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_17_LC_8_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_17_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_17_LC_8_21_3 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_17_LC_8_21_3  (
            .in0(N__29018),
            .in1(N__23450),
            .in2(N__23396),
            .in3(N__24698),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_8_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_8_21_4 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_8_21_4  (
            .in0(N__26763),
            .in1(N__23393),
            .in2(N__23384),
            .in3(N__23381),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(\delay_measurement_inst.un1_elapsed_time_hc_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_3_LC_8_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_3_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_3_LC_8_21_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_3_LC_8_21_5  (
            .in0(_gnd_net_),
            .in1(N__32790),
            .in2(N__23375),
            .in3(N__24240),
            .lcout(\delay_measurement_inst.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_22_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_22_0 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_22_0  (
            .in0(N__24221),
            .in1(_gnd_net_),
            .in2(N__30486),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_17_LC_8_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_17_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_17_LC_8_22_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_17_LC_8_22_1  (
            .in0(N__24550),
            .in1(N__28981),
            .in2(N__23462),
            .in3(N__23459),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_8_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_8_22_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_8_22_4  (
            .in0(N__30422),
            .in1(N__24485),
            .in2(_gnd_net_),
            .in3(N__33259),
            .lcout(),
            .ltout(\delay_measurement_inst.N_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_8_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_8_22_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_8_22_5 .LUT_INIT=16'b1111000011110101;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_8_22_5  (
            .in0(N__33130),
            .in1(_gnd_net_),
            .in2(N__23444),
            .in3(N__33378),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48354),
            .ce(),
            .sr(N__47878));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_8_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_8_22_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_8_22_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_8_22_6  (
            .in0(N__33377),
            .in1(N__33260),
            .in2(N__29207),
            .in3(N__33129),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48354),
            .ce(),
            .sr(N__47878));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_13_LC_8_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_13_LC_8_23_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_13_LC_8_23_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_13_LC_8_23_3  (
            .in0(N__34466),
            .in1(N__24308),
            .in2(_gnd_net_),
            .in3(N__33262),
            .lcout(\delay_measurement_inst.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_23_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_23_4  (
            .in0(N__29237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_23_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_23_5  (
            .in0(_gnd_net_),
            .in1(N__29271),
            .in2(_gnd_net_),
            .in3(N__29236),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_302_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_12_LC_8_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_12_LC_8_23_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_12_LC_8_23_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_12_LC_8_23_7  (
            .in0(N__33728),
            .in1(N__24341),
            .in2(_gnd_net_),
            .in3(N__33261),
            .lcout(\delay_measurement_inst.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_9_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_9_5_2 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_9_5_2  (
            .in0(N__24815),
            .in1(N__24831),
            .in2(_gnd_net_),
            .in3(N__30563),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48465),
            .ce(N__35904),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_9_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_9_6_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_9_6_1  (
            .in0(N__24814),
            .in1(N__24832),
            .in2(N__47927),
            .in3(N__30569),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48455),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_9_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_9_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__37996),
            .in2(_gnd_net_),
            .in3(N__23590),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_7_5  (
            .in0(N__27560),
            .in1(N__27401),
            .in2(N__29522),
            .in3(N__31912),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__23564),
            .in2(_gnd_net_),
            .in3(N__23542),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_8_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_8_0  (
            .in0(N__31512),
            .in1(N__29819),
            .in2(N__23515),
            .in3(N__26966),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_8_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__23507),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_9_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_9_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_9_8_2  (
            .in0(N__23702),
            .in1(N__27301),
            .in2(N__24884),
            .in3(N__24925),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_9_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_9_8_3 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_9_8_3  (
            .in0(N__24964),
            .in1(N__23648),
            .in2(N__23483),
            .in3(N__24728),
            .lcout(\current_shift_inst.PI_CTRL.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_9_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_9_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_9_8_4  (
            .in0(N__28463),
            .in1(N__31177),
            .in2(N__27776),
            .in3(N__31260),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_9_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_9_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_9_8_5  (
            .in0(N__24926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23742),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_8_7  (
            .in0(N__25016),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_9_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_9_0  (
            .in0(N__31517),
            .in1(N__29692),
            .in2(N__23655),
            .in3(N__27113),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23644),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_9_2 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_9_9_2  (
            .in0(N__27915),
            .in1(N__28282),
            .in2(N__28130),
            .in3(N__25100),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48427),
            .ce(),
            .sr(N__47796));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_9_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_9_9_3 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_9_9_3  (
            .in0(N__28279),
            .in1(N__28084),
            .in2(N__27965),
            .in3(N__25352),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48427),
            .ce(),
            .sr(N__47796));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_9_4 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_9_9_4  (
            .in0(N__28083),
            .in1(N__28280),
            .in2(N__27964),
            .in3(N__25325),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48427),
            .ce(),
            .sr(N__47796));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_9_6 .LUT_INIT=16'b0101111101010100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_9_9_6  (
            .in0(N__25283),
            .in1(N__28281),
            .in2(N__28131),
            .in3(N__27922),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48427),
            .ce(),
            .sr(N__47796));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_9_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_9_10_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__29906),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29933),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_10_2 .LUT_INIT=16'b0100010011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_9_10_2  (
            .in0(N__28122),
            .in1(N__27971),
            .in2(N__28304),
            .in3(N__25730),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_9_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_9_10_3 .LUT_INIT=16'b0101010100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_9_10_3  (
            .in0(N__25070),
            .in1(N__28285),
            .in2(N__28000),
            .in3(N__28125),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_9_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_9_10_4 .LUT_INIT=16'b0100010011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_9_10_4  (
            .in0(N__28121),
            .in1(N__27970),
            .in2(N__28303),
            .in3(N__25370),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_10_5 .LUT_INIT=16'b0000111110101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_9_10_5  (
            .in0(N__27969),
            .in1(N__28284),
            .in2(N__25580),
            .in3(N__28124),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_10_7 .LUT_INIT=16'b0000111110101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_9_10_7  (
            .in0(N__27968),
            .in1(N__28283),
            .in2(N__25295),
            .in3(N__28123),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(N__47799));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_9_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_9_11_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_9_11_0  (
            .in0(N__31469),
            .in1(N__30043),
            .in2(N__23703),
            .in3(N__27080),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_9_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_9_11_2 .LUT_INIT=16'b0000000111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_9_11_2  (
            .in0(N__28251),
            .in1(N__28129),
            .in2(N__28003),
            .in3(N__25037),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(N__47803));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_9_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_9_11_4 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_9_11_4  (
            .in0(N__28249),
            .in1(N__28127),
            .in2(N__28001),
            .in3(N__25607),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(N__47803));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_9_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_9_11_6 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_9_11_6  (
            .in0(N__28250),
            .in1(N__28128),
            .in2(N__28002),
            .in3(N__25550),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(N__47803));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_11_7 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_9_11_7  (
            .in0(N__28126),
            .in1(N__27981),
            .in2(N__25526),
            .in3(N__28252),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(N__47803));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_9_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_9_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_9_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29885),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_9_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_9_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_9_12_1 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_9_12_1  (
            .in0(N__28147),
            .in1(N__27985),
            .in2(N__25640),
            .in3(N__28247),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_12_2 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_9_12_2  (
            .in0(N__25229),
            .in1(_gnd_net_),
            .in2(N__28292),
            .in3(N__28152),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_3 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_3  (
            .in0(N__28148),
            .in1(N__27986),
            .in2(N__25514),
            .in3(N__28248),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_9_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_9_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_9_12_4 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_9_12_4  (
            .in0(N__28241),
            .in1(N__28150),
            .in2(N__28004),
            .in3(N__25499),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5  (
            .in0(N__28149),
            .in1(N__27987),
            .in2(N__25490),
            .in3(N__28246),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6  (
            .in0(N__28242),
            .in1(N__28151),
            .in2(N__28005),
            .in3(N__25478),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_9_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_9_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30047),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(N__47808));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_9_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_9_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_9_13_1  (
            .in0(N__27716),
            .in1(N__28712),
            .in2(N__27218),
            .in3(N__27629),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_9_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_9_13_2 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_9_13_2  (
            .in0(N__28253),
            .in1(N__28145),
            .in2(N__28006),
            .in3(N__25679),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48396),
            .ce(),
            .sr(N__47814));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28711),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_13_4 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_9_13_4  (
            .in0(N__28254),
            .in1(N__28146),
            .in2(N__28007),
            .in3(N__25661),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48396),
            .ce(),
            .sr(N__47814));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_13_5  (
            .in0(N__27208),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__23888),
            .in2(N__23876),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__23852),
            .in2(_gnd_net_),
            .in3(N__23834),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__23831),
            .in2(N__25760),
            .in3(N__23813),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23810),
            .in3(N__23789),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__23786),
            .in2(_gnd_net_),
            .in3(N__23768),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__24062),
            .in2(_gnd_net_),
            .in3(N__24044),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__24041),
            .in2(_gnd_net_),
            .in3(N__24023),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__24019),
            .in2(_gnd_net_),
            .in3(N__23999),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__23995),
            .in2(_gnd_net_),
            .in3(N__23975),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__23972),
            .in2(_gnd_net_),
            .in3(N__23954),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__23951),
            .in2(_gnd_net_),
            .in3(N__23933),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__23930),
            .in2(_gnd_net_),
            .in3(N__23912),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__23909),
            .in2(_gnd_net_),
            .in3(N__23891),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__24188),
            .in2(_gnd_net_),
            .in3(N__24170),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__24167),
            .in2(_gnd_net_),
            .in3(N__24149),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__25939),
            .in2(_gnd_net_),
            .in3(N__24146),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__24142),
            .in2(_gnd_net_),
            .in3(N__24122),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__24118),
            .in2(_gnd_net_),
            .in3(N__24098),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__24094),
            .in2(_gnd_net_),
            .in3(N__24080),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_9_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_9_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_9_16_3  (
            .in0(N__30765),
            .in1(N__32927),
            .in2(N__30296),
            .in3(N__30238),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_LC_9_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_LC_9_16_4 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_LC_9_16_4  (
            .in0(N__34429),
            .in1(N__30357),
            .in2(N__24071),
            .in3(N__24260),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt30 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlt30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_LC_9_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_LC_9_16_5 .LUT_INIT=16'b0011000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__36206),
            .in2(N__24266),
            .in3(N__34303),
            .lcout(\phase_controller_inst1.stoper_hc.un1_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_9_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_9_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_9_17_5  (
            .in0(N__33750),
            .in1(N__33698),
            .in2(N__34502),
            .in3(N__33581),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_LC_9_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_LC_9_17_6 .LUT_INIT=16'b0101000011010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_LC_9_17_6  (
            .in0(N__33635),
            .in1(N__24248),
            .in2(N__24263),
            .in3(N__30314),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_9_17_7.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_9_17_7.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_9_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_9_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47922),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_17_LC_9_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_17_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_17_LC_9_18_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_17_LC_9_18_0  (
            .in0(N__30229),
            .in1(N__24551),
            .in2(_gnd_net_),
            .in3(N__33289),
            .lcout(\delay_measurement_inst.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_9_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_9_18_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__32666),
            .in2(_gnd_net_),
            .in3(N__32716),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_9_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_9_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_9_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__25855),
            .in2(N__25921),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_9_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_9_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25882),
            .in2(N__25832),
            .in3(N__24194),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_9_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__25856),
            .in2(N__26194),
            .in3(N__24191),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_9_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_9_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__25828),
            .in2(N__26164),
            .in3(N__24458),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_9_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__26137),
            .in2(N__26195),
            .in3(N__24431),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_9_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__26116),
            .in2(N__26165),
            .in3(N__24398),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_9_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_9_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__26138),
            .in2(N__26089),
            .in3(N__24395),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_9_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__26117),
            .in2(N__26056),
            .in3(N__24371),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48366),
            .ce(N__24599),
            .sr(N__47859));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_9_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_9_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__26093),
            .in2(N__26029),
            .in3(N__24344),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_9_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_9_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__26002),
            .in2(N__26063),
            .in3(N__24311),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_9_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_9_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__26428),
            .in2(N__26030),
            .in3(N__24290),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_9_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__26003),
            .in2(N__26407),
            .in3(N__24578),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_9_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_9_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__26429),
            .in2(N__26381),
            .in3(N__24575),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_9_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__26350),
            .in2(N__26408),
            .in3(N__24554),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_9_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_9_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__26377),
            .in2(N__26326),
            .in3(N__24527),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_9_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_9_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__26351),
            .in2(N__26290),
            .in3(N__24524),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48360),
            .ce(N__24598),
            .sr(N__47865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_9_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__26327),
            .in2(N__26263),
            .in3(N__24497),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_9_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__26236),
            .in2(N__26297),
            .in3(N__24494),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_9_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__26215),
            .in2(N__26264),
            .in3(N__24491),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_9_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__26237),
            .in2(N__26641),
            .in3(N__24488),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_9_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__26216),
            .in2(N__26615),
            .in3(N__24626),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_9_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__26584),
            .in2(N__26642),
            .in3(N__24623),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_9_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__26611),
            .in2(N__26557),
            .in3(N__24620),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_9_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_9_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__26585),
            .in2(N__26524),
            .in3(N__24617),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48355),
            .ce(N__24597),
            .sr(N__47871));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_9_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__26494),
            .in2(N__26561),
            .in3(N__24614),
            .lcout(\delay_measurement_inst.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48349),
            .ce(N__24596),
            .sr(N__47875));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_9_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__26467),
            .in2(N__26531),
            .in3(N__24611),
            .lcout(\delay_measurement_inst.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48349),
            .ce(N__24596),
            .sr(N__47875));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_9_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__26447),
            .in2(N__26498),
            .in3(N__24608),
            .lcout(\delay_measurement_inst.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48349),
            .ce(N__24596),
            .sr(N__47875));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_9_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__26468),
            .in2(N__26783),
            .in3(N__24605),
            .lcout(\delay_measurement_inst.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48349),
            .ce(N__24596),
            .sr(N__47875));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_9_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_9_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24602),
            .lcout(\delay_measurement_inst.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48349),
            .ce(N__24596),
            .sr(N__47875));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_9_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_9_23_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_9_23_0  (
            .in0(N__26668),
            .in1(N__24688),
            .in2(N__29119),
            .in3(N__30640),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUV512_20_LC_9_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUV512_20_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUV512_20_LC_9_23_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUV512_20_LC_9_23_1  (
            .in0(N__29035),
            .in1(N__33376),
            .in2(N__24701),
            .in3(N__26702),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_28_LC_9_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_28_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_28_LC_9_23_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_28_LC_9_23_4  (
            .in0(N__29137),
            .in1(N__24689),
            .in2(_gnd_net_),
            .in3(N__33316),
            .lcout(\delay_measurement_inst.N_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_9_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_9_24_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_9_24_6  (
            .in0(N__24680),
            .in1(N__33437),
            .in2(_gnd_net_),
            .in3(N__33143),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48340),
            .ce(),
            .sr(N__47881));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6 (
            .in0(N__24674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_4_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_4_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_10_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24656),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48457),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24644),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_5_6  (
            .in0(N__43381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43419),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_5_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_5_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_5_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_5_7 (
            .in0(_gnd_net_),
            .in1(N__24632),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_10_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_10_6_0 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_10_6_0  (
            .in0(N__24813),
            .in1(N__24833),
            .in2(_gnd_net_),
            .in3(N__30564),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48437),
            .ce(),
            .sr(N__47774));
    defparam \delay_measurement_inst.prev_hc_sig_LC_10_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_10_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_10_6_1  (
            .in0(N__30565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48437),
            .ce(),
            .sr(N__47774));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36013),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48429),
            .ce(),
            .sr(N__47778));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_10_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_10_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29740),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48429),
            .ce(),
            .sr(N__47778));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_8_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_8_0  (
            .in0(N__31521),
            .in1(N__29771),
            .in2(N__24771),
            .in3(N__27140),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24761),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_10_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_10_8_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_10_8_2  (
            .in0(N__28299),
            .in1(N__28101),
            .in2(_gnd_net_),
            .in3(N__25160),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48419),
            .ce(),
            .sr(N__47784));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_8_4 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_10_8_4  (
            .in0(N__28300),
            .in1(N__28102),
            .in2(_gnd_net_),
            .in3(N__25127),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48419),
            .ce(),
            .sr(N__47784));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_10_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_10_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24727),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_8_7 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_8_7  (
            .in0(N__27131),
            .in1(N__29741),
            .in2(N__24744),
            .in3(N__31522),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_0 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_0  (
            .in0(N__26975),
            .in1(N__29861),
            .in2(N__25256),
            .in3(N__31514),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_9_1 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_9_1  (
            .in0(N__31547),
            .in1(N__31519),
            .in2(N__25028),
            .in3(N__27044),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_10_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_10_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31513),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_9_3 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_9_3  (
            .in0(N__29651),
            .in1(N__31520),
            .in2(N__31916),
            .in3(N__27170),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_4 .LUT_INIT=16'b0110011011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_4  (
            .in0(N__27065),
            .in1(N__29609),
            .in2(N__24980),
            .in3(N__31516),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_10_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_10_9_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_10_9_5  (
            .in0(N__31515),
            .in1(N__30014),
            .in2(N__24933),
            .in3(N__27092),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_10_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_10_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31735),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_9_7 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_9_7  (
            .in0(N__29630),
            .in1(N__31518),
            .in2(N__24893),
            .in3(N__27053),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__24844),
            .in2(N__24848),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_10_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__25252),
            .in2(N__25238),
            .in3(N__25220),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_10_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__25217),
            .in2(N__25208),
            .in3(N__25184),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_10_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__25181),
            .in2(N__25172),
            .in3(N__25151),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_10_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__25148),
            .in2(N__25139),
            .in3(N__25118),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__25115),
            .in2(N__25109),
            .in3(N__25094),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__25091),
            .in2(N__25085),
            .in3(N__25061),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__25769),
            .in2(N__27323),
            .in3(N__25058),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__25055),
            .in2(N__25049),
            .in3(N__25031),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__25472),
            .in2(N__25463),
            .in3(N__25436),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__25433),
            .in2(N__25424),
            .in3(N__25397),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__25394),
            .in2(N__25385),
            .in3(N__25364),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__25361),
            .in2(N__31868),
            .in3(N__25343),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__31556),
            .in2(N__25340),
            .in3(N__25313),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__31217),
            .in2(N__25310),
            .in3(N__25286),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__31133),
            .in2(N__29666),
            .in3(N__25274),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__27350),
            .in2(N__25271),
            .in3(N__25628),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__28412),
            .in2(N__25625),
            .in3(N__25601),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__27509),
            .in2(N__25598),
            .in3(N__25568),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__29540),
            .in2(N__25565),
            .in3(N__25544),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__27467),
            .in2(N__25541),
            .in3(N__25517),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__27485),
            .in2(N__29465),
            .in3(N__25502),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__27338),
            .in2(N__26954),
            .in3(N__25493),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(N__27497),
            .in2(N__30953),
            .in3(N__25481),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__27413),
            .in2(N__25799),
            .in3(N__25751),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__27671),
            .in2(N__25748),
            .in3(N__25721),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__27596),
            .in2(N__25718),
            .in3(N__25691),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__28688),
            .in2(N__25688),
            .in3(N__25673),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__27182),
            .in2(N__25670),
            .in3(N__25655),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__25790),
            .in2(N__28681),
            .in3(N__25652),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__28677),
            .in2(N__25778),
            .in3(N__25649),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__25784),
            .in2(N__28682),
            .in3(N__25646),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_14_0  (
            .in0(N__27879),
            .in1(N__31523),
            .in2(_gnd_net_),
            .in3(N__25643),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27453),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_10_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28374),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27747),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_10_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_10_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28326),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27275),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__25974),
            .in2(_gnd_net_),
            .in3(N__35619),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_15_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_15_2  (
            .in0(N__35502),
            .in1(N__35289),
            .in2(_gnd_net_),
            .in3(N__35377),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_10_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_10_15_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_10_15_7  (
            .in0(N__45523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45482),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__34612),
            .in2(_gnd_net_),
            .in3(N__33798),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_10_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_16_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_10_16_1  (
            .in0(N__35491),
            .in1(N__28880),
            .in2(N__25982),
            .in3(N__45488),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48372),
            .ce(),
            .sr(N__47820));
    defparam \phase_controller_inst1.state_2_LC_10_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_10_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_10_16_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_10_16_3  (
            .in0(N__33799),
            .in1(N__30703),
            .in2(N__34616),
            .in3(N__30678),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48372),
            .ce(),
            .sr(N__47820));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_16_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__35288),
            .in2(_gnd_net_),
            .in3(N__35376),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_16_5 .LUT_INIT=16'b1100100011011000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_10_16_5  (
            .in0(N__25955),
            .in1(N__30679),
            .in2(N__25949),
            .in3(N__35631),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48372),
            .ce(),
            .sr(N__47820));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_16_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_16_6  (
            .in0(N__35290),
            .in1(N__35492),
            .in2(N__35422),
            .in3(N__25946),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48372),
            .ce(),
            .sr(N__47820));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_10_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_10_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_10_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_10_17_0  (
            .in0(N__26936),
            .in1(N__25908),
            .in2(_gnd_net_),
            .in3(N__25892),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_10_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_10_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_10_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_10_17_1  (
            .in0(N__26932),
            .in1(N__25875),
            .in2(_gnd_net_),
            .in3(N__25859),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_10_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_10_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_10_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_10_17_2  (
            .in0(N__26937),
            .in1(N__25854),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_10_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_10_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_10_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_10_17_3  (
            .in0(N__26933),
            .in1(N__25824),
            .in2(_gnd_net_),
            .in3(N__25802),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_10_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_10_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_10_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_10_17_4  (
            .in0(N__26938),
            .in1(N__26182),
            .in2(_gnd_net_),
            .in3(N__26168),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_10_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_10_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_10_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_10_17_5  (
            .in0(N__26934),
            .in1(N__26157),
            .in2(_gnd_net_),
            .in3(N__26141),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_10_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_10_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_10_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_10_17_6  (
            .in0(N__26939),
            .in1(N__26136),
            .in2(_gnd_net_),
            .in3(N__26120),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_10_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_10_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_10_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_10_17_7  (
            .in0(N__26935),
            .in1(N__26110),
            .in2(_gnd_net_),
            .in3(N__26096),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__48367),
            .ce(N__28948),
            .sr(N__47827));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_10_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_10_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_10_18_0  (
            .in0(N__26927),
            .in1(N__26085),
            .in2(_gnd_net_),
            .in3(N__26066),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_10_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_10_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_10_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_10_18_1  (
            .in0(N__26931),
            .in1(N__26055),
            .in2(_gnd_net_),
            .in3(N__26033),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_10_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_10_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_10_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_10_18_2  (
            .in0(N__26924),
            .in1(N__26022),
            .in2(_gnd_net_),
            .in3(N__26006),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_10_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_10_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_10_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_10_18_3  (
            .in0(N__26928),
            .in1(N__26001),
            .in2(_gnd_net_),
            .in3(N__25985),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_10_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_10_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_10_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_10_18_4  (
            .in0(N__26925),
            .in1(N__26427),
            .in2(_gnd_net_),
            .in3(N__26411),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_10_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_10_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_10_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_10_18_5  (
            .in0(N__26929),
            .in1(N__26400),
            .in2(_gnd_net_),
            .in3(N__26384),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_10_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_10_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_10_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_10_18_6  (
            .in0(N__26926),
            .in1(N__26373),
            .in2(_gnd_net_),
            .in3(N__26354),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_10_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_10_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_10_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_10_18_7  (
            .in0(N__26930),
            .in1(N__26344),
            .in2(_gnd_net_),
            .in3(N__26330),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__48362),
            .ce(N__28949),
            .sr(N__47836));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_10_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_10_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_10_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_10_19_0  (
            .in0(N__26910),
            .in1(N__26322),
            .in2(_gnd_net_),
            .in3(N__26300),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_10_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_10_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_10_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_10_19_1  (
            .in0(N__26917),
            .in1(N__26289),
            .in2(_gnd_net_),
            .in3(N__26267),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_10_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_10_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_10_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_10_19_2  (
            .in0(N__26911),
            .in1(N__26256),
            .in2(_gnd_net_),
            .in3(N__26240),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_10_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_10_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_10_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_10_19_3  (
            .in0(N__26914),
            .in1(N__26235),
            .in2(_gnd_net_),
            .in3(N__26219),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_10_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_10_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_10_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_10_19_4  (
            .in0(N__26912),
            .in1(N__26214),
            .in2(_gnd_net_),
            .in3(N__26198),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_10_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_10_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_10_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_10_19_5  (
            .in0(N__26915),
            .in1(N__26634),
            .in2(_gnd_net_),
            .in3(N__26618),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_10_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_10_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_10_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_10_19_6  (
            .in0(N__26913),
            .in1(N__26607),
            .in2(_gnd_net_),
            .in3(N__26588),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_10_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_10_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_10_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_10_19_7  (
            .in0(N__26916),
            .in1(N__26578),
            .in2(_gnd_net_),
            .in3(N__26564),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__48356),
            .ce(N__28940),
            .sr(N__47847));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_10_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_10_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_10_20_0  (
            .in0(N__26918),
            .in1(N__26553),
            .in2(_gnd_net_),
            .in3(N__26534),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__48350),
            .ce(N__28944),
            .sr(N__47852));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_10_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_10_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_10_20_1  (
            .in0(N__26922),
            .in1(N__26523),
            .in2(_gnd_net_),
            .in3(N__26501),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__48350),
            .ce(N__28944),
            .sr(N__47852));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_10_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_10_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_10_20_2  (
            .in0(N__26919),
            .in1(N__26487),
            .in2(_gnd_net_),
            .in3(N__26471),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__48350),
            .ce(N__28944),
            .sr(N__47852));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_10_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_10_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_10_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_10_20_3  (
            .in0(N__26923),
            .in1(N__26466),
            .in2(_gnd_net_),
            .in3(N__26450),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__48350),
            .ce(N__28944),
            .sr(N__47852));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_10_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_10_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_10_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_10_20_4  (
            .in0(N__26920),
            .in1(N__26446),
            .in2(_gnd_net_),
            .in3(N__26432),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__48350),
            .ce(N__28944),
            .sr(N__47852));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_10_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_10_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_10_20_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_10_20_5  (
            .in0(N__26779),
            .in1(N__26921),
            .in2(_gnd_net_),
            .in3(N__26786),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48350),
            .ce(N__28944),
            .sr(N__47852));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_15_LC_10_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_15_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_15_LC_10_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_15_LC_10_21_3  (
            .in0(N__34400),
            .in1(N__26765),
            .in2(_gnd_net_),
            .in3(N__33293),
            .lcout(),
            .ltout(\delay_measurement_inst.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_10_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_10_21_4 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__33414),
            .in2(N__26744),
            .in3(N__33077),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48346),
            .ce(),
            .sr(N__47860));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_10_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_10_21_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_10_21_5  (
            .in0(N__26741),
            .in1(N__26735),
            .in2(N__26729),
            .in3(N__26720),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_10_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_10_22_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__26714),
            .in2(_gnd_net_),
            .in3(N__26708),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI45SG1_21_LC_10_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI45SG1_21_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI45SG1_21_LC_10_22_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI45SG1_21_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26696),
            .in3(N__26693),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_1_LC_10_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_1_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_1_LC_10_22_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_1_LC_10_22_5  (
            .in0(N__32866),
            .in1(N__33315),
            .in2(_gnd_net_),
            .in3(N__26687),
            .lcout(\delay_measurement_inst.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_27_LC_10_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_27_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_27_LC_10_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_27_LC_10_23_6  (
            .in0(N__26669),
            .in1(N__29096),
            .in2(_gnd_net_),
            .in3(N__33317),
            .lcout(\delay_measurement_inst.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_10_27_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_10_27_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_10_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35831),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48330),
            .ce(),
            .sr(N__47884));
    defparam \delay_measurement_inst.tr_state_0_LC_11_3_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_11_3_5 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_11_3_5  (
            .in0(N__29366),
            .in1(N__29343),
            .in2(_gnd_net_),
            .in3(N__29327),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48458),
            .ce(N__35927),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_4_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_4_6  (
            .in0(N__39072),
            .in1(N__39114),
            .in2(N__38748),
            .in3(N__42747),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_11_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_11_5_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_11_5_0  (
            .in0(N__41433),
            .in1(N__41288),
            .in2(_gnd_net_),
            .in3(N__37276),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48438),
            .ce(N__30869),
            .sr(N__47765));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_5_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_5_1  (
            .in0(N__29414),
            .in1(N__41429),
            .in2(_gnd_net_),
            .in3(N__40985),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48438),
            .ce(N__30869),
            .sr(N__47765));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_5_2 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_5_2  (
            .in0(N__40880),
            .in1(_gnd_net_),
            .in2(N__41435),
            .in3(N__37275),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48438),
            .ce(N__30869),
            .sr(N__47765));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_5_3 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_5_3  (
            .in0(N__37277),
            .in1(N__41434),
            .in2(_gnd_net_),
            .in3(N__41234),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48438),
            .ce(N__30869),
            .sr(N__47765));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31854),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_11_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_11_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_11_6_3  (
            .in0(N__39063),
            .in1(N__39113),
            .in2(N__38747),
            .in3(N__42746),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_11_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_11_6_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_11_6_6  (
            .in0(N__40936),
            .in1(N__41128),
            .in2(N__30890),
            .in3(N__37261),
            .lcout(\delay_measurement_inst.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_11_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_11_6_7 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_11_6_7  (
            .in0(N__37262),
            .in1(N__40937),
            .in2(N__40835),
            .in3(N__40984),
            .lcout(\delay_measurement_inst.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_11_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_11_7_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_11_7_0  (
            .in0(N__37582),
            .in1(N__45487),
            .in2(N__28789),
            .in3(N__27038),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48420),
            .ce(),
            .sr(N__47775));
    defparam \phase_controller_inst1.start_timer_tr_LC_11_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_7_5 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_11_7_5  (
            .in0(N__45486),
            .in1(N__43601),
            .in2(N__27029),
            .in3(N__43855),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48420),
            .ce(),
            .sr(N__47775));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__26999),
            .in2(_gnd_net_),
            .in3(N__27010),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__26993),
            .in2(_gnd_net_),
            .in3(N__29932),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__26987),
            .in2(_gnd_net_),
            .in3(N__29905),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__26981),
            .in2(_gnd_net_),
            .in3(N__29881),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__29588),
            .in2(_gnd_net_),
            .in3(N__26969),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__29432),
            .in2(_gnd_net_),
            .in3(N__26957),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__29582),
            .in2(_gnd_net_),
            .in3(N__27134),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__29426),
            .in2(_gnd_net_),
            .in3(N__27125),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__27122),
            .in2(_gnd_net_),
            .in3(N__27104),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__27101),
            .in2(_gnd_net_),
            .in3(N__27086),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29447),
            .in3(N__27083),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__29438),
            .in2(_gnd_net_),
            .in3(N__27068),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__29604),
            .in2(_gnd_net_),
            .in3(N__27056),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__29625),
            .in2(_gnd_net_),
            .in3(N__27047),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__31546),
            .in2(_gnd_net_),
            .in3(N__27173),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__29646),
            .in2(_gnd_net_),
            .in3(N__27164),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__31634),
            .in2(_gnd_net_),
            .in3(N__27161),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__31298),
            .in2(_gnd_net_),
            .in3(N__27158),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__31205),
            .in2(_gnd_net_),
            .in3(N__27155),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__31117),
            .in2(_gnd_net_),
            .in3(N__27152),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__31063),
            .in2(_gnd_net_),
            .in3(N__27149),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__28574),
            .in2(_gnd_net_),
            .in3(N__27146),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__29569),
            .in2(_gnd_net_),
            .in3(N__27143),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__28522),
            .in2(_gnd_net_),
            .in3(N__27251),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__31093),
            .in2(_gnd_net_),
            .in3(N__27248),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__28546),
            .in2(_gnd_net_),
            .in3(N__27245),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__31042),
            .in2(_gnd_net_),
            .in3(N__27242),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__28498),
            .in2(_gnd_net_),
            .in3(N__27239),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__28900),
            .in2(_gnd_net_),
            .in3(N__27236),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__27665),
            .in2(_gnd_net_),
            .in3(N__27233),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__27590),
            .in2(_gnd_net_),
            .in3(N__27230),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_11_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_11_7  (
            .in0(N__31428),
            .in1(N__27227),
            .in2(_gnd_net_),
            .in3(N__27185),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_11_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_11_12_0 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_11_12_0  (
            .in0(N__28573),
            .in1(N__31422),
            .in2(N__27575),
            .in3(N__27518),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_12_1 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_12_1  (
            .in0(N__31426),
            .in1(N__31043),
            .in2(N__31684),
            .in3(N__27503),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_11_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_11_12_3 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_11_12_3  (
            .in0(N__31424),
            .in1(N__27491),
            .in2(N__29517),
            .in3(N__31094),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_11_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_11_12_4 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_11_12_4  (
            .in0(N__28523),
            .in1(N__31795),
            .in2(N__27479),
            .in3(N__31423),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_11_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_11_12_5 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_11_12_5  (
            .in0(N__31427),
            .in1(N__27457),
            .in2(N__28499),
            .in3(N__27419),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_11_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_11_12_6 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_11_12_6  (
            .in0(N__31121),
            .in1(N__31421),
            .in2(N__27407),
            .in3(N__27359),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_12_7 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_12_7  (
            .in0(N__31425),
            .in1(N__28547),
            .in2(N__31856),
            .in3(N__27344),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_13_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_13_0  (
            .in0(N__29972),
            .in1(N__31511),
            .in2(N__27293),
            .in3(N__27332),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_11_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_11_13_2 .LUT_INIT=16'b0000000111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_11_13_2  (
            .in0(N__28295),
            .in1(N__28157),
            .in2(N__27884),
            .in3(N__27311),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48384),
            .ce(),
            .sr(N__47800));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_13_3 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_11_13_3  (
            .in0(N__28153),
            .in1(N__28296),
            .in2(N__27880),
            .in3(N__28403),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48384),
            .ce(),
            .sr(N__47800));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_13_4 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_11_13_4  (
            .in0(N__28293),
            .in1(N__28155),
            .in2(N__27882),
            .in3(N__28358),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48384),
            .ce(),
            .sr(N__47800));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_11_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_11_13_5 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_11_13_5  (
            .in0(N__28154),
            .in1(N__28297),
            .in2(N__27881),
            .in3(N__28310),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48384),
            .ce(),
            .sr(N__47800));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_11_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_11_13_6 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_11_13_6  (
            .in0(N__28294),
            .in1(N__28156),
            .in2(N__27883),
            .in3(N__27782),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48384),
            .ce(),
            .sr(N__47800));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_11_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_11_14_0 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_11_14_0  (
            .in0(N__31506),
            .in1(N__28901),
            .in2(N__27731),
            .in3(N__27680),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_11_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_11_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__27664),
            .in2(_gnd_net_),
            .in3(N__31504),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_11_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_11_14_2 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_11_14_2  (
            .in0(N__31507),
            .in1(N__27650),
            .in2(N__27608),
            .in3(N__27605),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_11_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_11_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_11_14_3  (
            .in0(N__27589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31505),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_11_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_11_14_4 .LUT_INIT=16'b0111110101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_11_14_4  (
            .in0(N__31508),
            .in1(N__28742),
            .in2(N__28733),
            .in3(N__28730),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_11_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_11_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31509),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_11_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_11_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_11_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_11_14_6  (
            .in0(N__31510),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48378),
            .ce(),
            .sr(N__47804));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__28569),
            .in2(_gnd_net_),
            .in3(N__31497),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_15_1  (
            .in0(N__31500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28545),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_15_2  (
            .in0(N__29568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31498),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_3  (
            .in0(N__31499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28515),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_15_4  (
            .in0(N__28491),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31501),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_11_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_11_15_5 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_11_15_5  (
            .in0(N__31503),
            .in1(N__31070),
            .in2(N__28472),
            .in3(N__28424),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_11_15_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_11_15_6  (
            .in0(N__36606),
            .in1(N__36471),
            .in2(_gnd_net_),
            .in3(N__36323),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_15_7  (
            .in0(N__31502),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28899),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__30702),
            .in2(_gnd_net_),
            .in3(N__30677),
            .lcout(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_2 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_2  (
            .in0(N__36208),
            .in1(N__36148),
            .in2(_gnd_net_),
            .in3(N__36122),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48363),
            .ce(N__28843),
            .sr(N__47821));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_17_3 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_11_17_3  (
            .in0(N__32935),
            .in1(N__33957),
            .in2(_gnd_net_),
            .in3(N__34270),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48363),
            .ce(N__28843),
            .sr(N__47821));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_11_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_11_18_0 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_11_18_0  (
            .in0(N__33090),
            .in1(N__33499),
            .in2(N__30509),
            .in3(N__33325),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48357),
            .ce(),
            .sr(N__47828));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_11_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_11_18_1 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_11_18_1  (
            .in0(N__33324),
            .in1(N__32565),
            .in2(N__33522),
            .in3(N__33089),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48357),
            .ce(),
            .sr(N__47828));
    defparam \phase_controller_inst2.state_3_LC_11_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_11_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_11_18_4 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.state_3_LC_11_18_4  (
            .in0(N__35789),
            .in1(N__28793),
            .in2(N__35822),
            .in3(N__33769),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48357),
            .ce(),
            .sr(N__47828));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_9_LC_11_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_9_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_9_LC_11_19_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_9_LC_11_19_0  (
            .in0(N__33619),
            .in1(N__28763),
            .in2(_gnd_net_),
            .in3(N__33321),
            .lcout(),
            .ltout(\delay_measurement_inst.N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_11_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_11_19_1 .LUT_INIT=16'b1111000011110101;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_11_19_1  (
            .in0(N__33513),
            .in1(_gnd_net_),
            .in2(N__29069),
            .in3(N__33076),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48351),
            .ce(),
            .sr(N__47837));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_11_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_11_19_3 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_11_19_3  (
            .in0(N__33512),
            .in1(N__29066),
            .in2(_gnd_net_),
            .in3(N__33075),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48351),
            .ce(),
            .sr(N__47837));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_2_LC_11_20_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_2_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_2_LC_11_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_2_LC_11_20_2  (
            .in0(N__33313),
            .in1(N__34039),
            .in2(_gnd_net_),
            .in3(N__29057),
            .lcout(\delay_measurement_inst.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46379_20_LC_11_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46379_20_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46379_20_LC_11_20_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46379_20_LC_11_20_3  (
            .in0(N__29039),
            .in1(N__29017),
            .in2(N__29003),
            .in3(N__28991),
            .lcout(\delay_measurement_inst.delay_hc_reg3lt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_18_LC_11_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_18_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_18_LC_11_20_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_18_LC_11_20_5  (
            .in0(N__30748),
            .in1(N__28982),
            .in2(_gnd_net_),
            .in3(N__33312),
            .lcout(\delay_measurement_inst.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_20_7 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_20_7  (
            .in0(N__29305),
            .in1(N__29278),
            .in2(_gnd_net_),
            .in3(N__29226),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_303_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_11_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_11_21_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_11_21_0  (
            .in0(N__33475),
            .in1(N__33308),
            .in2(N__29189),
            .in3(N__33042),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48342),
            .ce(),
            .sr(N__47853));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_11_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_11_21_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_11_21_1  (
            .in0(N__33045),
            .in1(N__33478),
            .in2(_gnd_net_),
            .in3(N__28910),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48342),
            .ce(),
            .sr(N__47853));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_11_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_11_21_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_11_21_2  (
            .in0(N__33477),
            .in1(N__30629),
            .in2(_gnd_net_),
            .in3(N__33044),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48342),
            .ce(),
            .sr(N__47853));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_11_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_11_21_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_11_21_3  (
            .in0(N__29309),
            .in1(N__29282),
            .in2(_gnd_net_),
            .in3(N__29227),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48342),
            .ce(),
            .sr(N__47853));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_11_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_11_21_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_11_21_6  (
            .in0(N__33474),
            .in1(N__33307),
            .in2(N__29156),
            .in3(N__33041),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48342),
            .ce(),
            .sr(N__47853));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_11_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_11_21_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_11_21_7 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_11_21_7  (
            .in0(N__33043),
            .in1(N__29170),
            .in2(N__33326),
            .in3(N__33476),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48342),
            .ce(),
            .sr(N__47853));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_11_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_11_22_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_11_22_0  (
            .in0(N__29203),
            .in1(N__29185),
            .in2(N__29174),
            .in3(N__29152),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_11_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_11_22_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_11_22_1  (
            .in0(N__29141),
            .in1(N__29092),
            .in2(N__29123),
            .in3(N__30611),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_30_LC_11_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_30_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_30_LC_11_22_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_30_LC_11_22_7  (
            .in0(N__30599),
            .in1(N__29120),
            .in2(_gnd_net_),
            .in3(N__33320),
            .lcout(\delay_measurement_inst.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_11_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_11_23_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_11_23_0  (
            .in0(N__33511),
            .in1(N__29102),
            .in2(_gnd_net_),
            .in3(N__33123),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48336),
            .ce(),
            .sr(N__47866));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_11_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_11_23_2 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_11_23_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_11_23_2  (
            .in0(N__33510),
            .in1(N__29081),
            .in2(_gnd_net_),
            .in3(N__33122),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48336),
            .ce(),
            .sr(N__47866));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_1_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_1_1  (
            .in0(_gnd_net_),
            .in1(N__42606),
            .in2(_gnd_net_),
            .in3(N__42582),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_304_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_2_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_2_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_12_2_1  (
            .in0(N__29363),
            .in1(N__29345),
            .in2(N__47926),
            .in3(N__29326),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48456),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR1_LC_12_2_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_12_2_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_12_2_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_12_2_5 (
            .in0(N__29384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48456),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_12_2_7.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_12_2_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_12_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_12_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29372),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48456),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_3_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29365),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48445),
            .ce(),
            .sr(N__47746));
    defparam \delay_measurement_inst.start_timer_tr_LC_12_3_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_3_7 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_12_3_7  (
            .in0(N__29364),
            .in1(N__29344),
            .in2(_gnd_net_),
            .in3(N__29325),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48445),
            .ce(),
            .sr(N__47746));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_4_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_4_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_4_2 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_12_4_2  (
            .in0(N__42634),
            .in1(N__42616),
            .in2(_gnd_net_),
            .in3(N__42581),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48436),
            .ce(),
            .sr(N__47752));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__47918),
            .in2(_gnd_net_),
            .in3(N__39277),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_12_5_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_12_5_6 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_12_5_6  (
            .in0(N__30938),
            .in1(N__40692),
            .in2(_gnd_net_),
            .in3(N__39250),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48428),
            .ce(N__30868),
            .sr(N__47757));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_5_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_5_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_5_7 .LUT_INIT=16'b1010111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_5_7  (
            .in0(N__39249),
            .in1(N__30937),
            .in2(N__40702),
            .in3(N__45649),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48428),
            .ce(N__30868),
            .sr(N__47757));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_12_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_12_6_0 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_12_6_0  (
            .in0(N__40701),
            .in1(N__45599),
            .in2(N__39260),
            .in3(N__30936),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_12_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_12_6_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_12_6_1  (
            .in0(N__29412),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__41008),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_12_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_12_6_2 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_12_6_2  (
            .in0(N__41129),
            .in1(N__29413),
            .in2(N__41427),
            .in3(N__29420),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_12_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_12_6_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_12_6_4  (
            .in0(N__41406),
            .in1(N__29409),
            .in2(_gnd_net_),
            .in3(N__41078),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_6_5 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_6_5  (
            .in0(N__41261),
            .in1(N__41410),
            .in2(_gnd_net_),
            .in3(N__37257),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_12_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_12_6_6 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_12_6_6  (
            .in0(N__41407),
            .in1(N__29410),
            .in2(_gnd_net_),
            .in3(N__41054),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_12_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_12_6_7 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_12_6_7  (
            .in0(N__29411),
            .in1(N__41408),
            .in2(_gnd_net_),
            .in3(N__41033),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(N__30870),
            .sr(N__47766));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_7_0  (
            .in0(N__41032),
            .in1(N__41053),
            .in2(N__41009),
            .in3(N__41074),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ),
            .ltout(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_7_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_7_1  (
            .in0(N__41149),
            .in1(N__40630),
            .in2(N__29390),
            .in3(N__37245),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_7_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29387),
            .in3(N__40924),
            .lcout(\delay_measurement_inst.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29518),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_7_5  (
            .in0(N__40975),
            .in1(N__41111),
            .in2(N__40934),
            .in3(N__40690),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_7_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_7_6  (
            .in0(N__37576),
            .in1(N__37511),
            .in2(_gnd_net_),
            .in3(N__37783),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_12_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_12_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__38549),
            .in2(_gnd_net_),
            .in3(N__38488),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48402),
            .ce(N__42683),
            .sr(N__47776));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_12_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_12_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__38067),
            .in2(_gnd_net_),
            .in3(N__39332),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48402),
            .ce(N__42683),
            .sr(N__47776));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29971),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30042),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29814),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29733),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_12_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_12_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31181),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_1  (
            .in0(N__31431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29650),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35972),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_12_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_12_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_12_9_3  (
            .in0(N__31430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29629),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_12_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_12_9_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__31429),
            .in2(_gnd_net_),
            .in3(N__29608),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29850),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29760),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_12_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_12_9_7 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_12_9_7  (
            .in0(N__31432),
            .in1(N__29576),
            .in2(N__31745),
            .in3(N__29546),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0  (
            .in0(N__36014),
            .in1(N__29528),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30200),
            .in3(N__29915),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__29912),
            .in2(_gnd_net_),
            .in3(N__29888),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__30305),
            .in2(_gnd_net_),
            .in3(N__29864),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__32255),
            .in2(_gnd_net_),
            .in3(N__29834),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__29831),
            .in2(_gnd_net_),
            .in3(N__29789),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__29786),
            .in2(_gnd_net_),
            .in3(N__29744),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__32267),
            .in2(_gnd_net_),
            .in3(N__29711),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__48392),
            .ce(),
            .sr(N__47785));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__29708),
            .in2(_gnd_net_),
            .in3(N__29669),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_8 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__30254),
            .in2(_gnd_net_),
            .in3(N__30053),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__36770),
            .in2(_gnd_net_),
            .in3(N__30050),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__30173),
            .in2(_gnd_net_),
            .in3(N__30020),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__36650),
            .in2(_gnd_net_),
            .in3(N__30017),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_12_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_12_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30006),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_11_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_11_7  (
            .in0(N__36477),
            .in1(N__36324),
            .in2(N__36629),
            .in3(N__30101),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48388),
            .ce(),
            .sr(N__47789));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_12_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_12_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29970),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_12_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_12_1  (
            .in0(N__36464),
            .in1(N__36619),
            .in2(N__30089),
            .in3(N__36328),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_12_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_12_2  (
            .in0(N__36325),
            .in1(N__36468),
            .in2(N__36626),
            .in3(N__30074),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_12_3 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_12_3  (
            .in0(N__36465),
            .in1(N__36620),
            .in2(N__30065),
            .in3(N__36329),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_12_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_12_4  (
            .in0(N__36326),
            .in1(N__36469),
            .in2(N__36627),
            .in3(N__30161),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_12_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_12_5  (
            .in0(N__36466),
            .in1(N__36621),
            .in2(N__30152),
            .in3(N__36330),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_12_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_12_6  (
            .in0(N__36327),
            .in1(N__36470),
            .in2(N__36628),
            .in3(N__30140),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_12_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_12_7  (
            .in0(N__36467),
            .in1(N__36622),
            .in2(N__30131),
            .in3(N__36331),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(N__47792));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__35705),
            .in2(N__35690),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_12_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_12_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__32105),
            .in2(_gnd_net_),
            .in3(N__30092),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_12_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_12_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__36026),
            .in2(N__32084),
            .in3(N__30077),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_12_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_12_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__32063),
            .in2(_gnd_net_),
            .in3(N__30068),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_12_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_12_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__32045),
            .in2(_gnd_net_),
            .in3(N__30056),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_12_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_12_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__32012),
            .in2(_gnd_net_),
            .in3(N__30155),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_12_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_12_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__31994),
            .in2(_gnd_net_),
            .in3(N__30143),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_12_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_12_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__31976),
            .in2(_gnd_net_),
            .in3(N__30134),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_12_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_12_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__31940),
            .in2(_gnd_net_),
            .in3(N__30119),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_12_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_12_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__35651),
            .in2(_gnd_net_),
            .in3(N__30116),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_12_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_12_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__35723),
            .in2(_gnd_net_),
            .in3(N__30113),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_12_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_12_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__32236),
            .in2(_gnd_net_),
            .in3(N__30110),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_12_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_12_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__32215),
            .in2(_gnd_net_),
            .in3(N__30107),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_12_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_12_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__32194),
            .in2(_gnd_net_),
            .in3(N__30104),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_12_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_12_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__32521),
            .in2(_gnd_net_),
            .in3(N__30188),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_12_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_12_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__32501),
            .in2(_gnd_net_),
            .in3(N__30185),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_12_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_12_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__32483),
            .in2(_gnd_net_),
            .in3(N__30182),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_12_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_12_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__32465),
            .in2(_gnd_net_),
            .in3(N__30179),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_12_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_12_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__32447),
            .in2(_gnd_net_),
            .in3(N__30176),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36646),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_12_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_12_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_12_16_0 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_12_16_0  (
            .in0(N__34129),
            .in1(N__33922),
            .in2(N__30361),
            .in3(N__34291),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48361),
            .ce(N__36076),
            .sr(N__47809));
    defparam \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_12_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_12_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_12_16_1 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_12_16_1  (
            .in0(N__34289),
            .in1(N__30447),
            .in2(N__33961),
            .in3(N__34128),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48361),
            .ce(N__36076),
            .sr(N__47809));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_12_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_12_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_12_16_2 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_12_16_2  (
            .in0(N__34130),
            .in1(N__33923),
            .in2(N__33644),
            .in3(N__34292),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48361),
            .ce(N__36076),
            .sr(N__47809));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_12_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_12_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_12_16_4 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_12_16_4  (
            .in0(N__30242),
            .in1(N__33921),
            .in2(_gnd_net_),
            .in3(N__34290),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48361),
            .ce(N__36076),
            .sr(N__47809));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_12_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_12_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_12_16_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_12_16_5  (
            .in0(N__34288),
            .in1(N__30766),
            .in2(_gnd_net_),
            .in3(N__33936),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48361),
            .ce(N__36076),
            .sr(N__47809));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_16_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_16_7  (
            .in0(N__34428),
            .in1(N__30353),
            .in2(N__32936),
            .in3(N__34507),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_12_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_12_17_1 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto6_LC_12_17_1  (
            .in0(N__32364),
            .in1(N__32430),
            .in2(N__30451),
            .in3(N__30515),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35951),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_12_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_12_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_12_17_6  (
            .in0(N__30505),
            .in1(N__32969),
            .in2(N__30392),
            .in3(N__30295),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36668),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_12_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_12_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_12_18_0  (
            .in0(N__32674),
            .in1(N__30231),
            .in2(N__30764),
            .in3(N__32725),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35987),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_18_2 .LUT_INIT=16'b0000110001001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_18_2  (
            .in0(N__34044),
            .in1(N__30398),
            .in2(N__32789),
            .in3(N__32871),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_12_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_12_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_12_18_3  (
            .in0(N__33533),
            .in1(N__30533),
            .in2(N__30527),
            .in3(N__30524),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_18_4  (
            .in0(N__34043),
            .in1(N__32558),
            .in2(N__32788),
            .in3(N__32870),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_12_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_12_18_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_12_18_7  (
            .in0(N__30504),
            .in1(N__32968),
            .in2(N__30387),
            .in3(N__36123),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_5_LC_12_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_5_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_5_LC_12_19_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_5_LC_12_19_4  (
            .in0(N__32357),
            .in1(N__30488),
            .in2(_gnd_net_),
            .in3(N__33322),
            .lcout(),
            .ltout(\delay_measurement_inst.N_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_12_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_12_19_5 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__33521),
            .in2(N__30455),
            .in3(N__33059),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48345),
            .ce(),
            .sr(N__47829));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_19_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_19_6  (
            .in0(N__30434),
            .in1(N__32356),
            .in2(_gnd_net_),
            .in3(N__32425),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_12_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_12_19_7 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_12_19_7  (
            .in0(N__33323),
            .in1(N__33520),
            .in2(N__30391),
            .in3(N__33058),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48345),
            .ce(),
            .sr(N__47829));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_12_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_12_20_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_12_20_0  (
            .in0(N__33516),
            .in1(N__33314),
            .in2(N__36205),
            .in3(N__33046),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48341),
            .ce(),
            .sr(N__47838));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_12_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_12_20_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_12_20_1  (
            .in0(N__33047),
            .in1(N__33517),
            .in2(_gnd_net_),
            .in3(N__30776),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48341),
            .ce(),
            .sr(N__47838));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_12_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_12_20_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_12_20_5  (
            .in0(N__33048),
            .in1(N__33518),
            .in2(_gnd_net_),
            .in3(N__30719),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48341),
            .ce(),
            .sr(N__47838));
    defparam \phase_controller_inst1.state_1_LC_12_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_20_6 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_20_6  (
            .in0(N__43442),
            .in1(N__30713),
            .in2(N__43367),
            .in3(N__30686),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48341),
            .ce(),
            .sr(N__47838));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_12_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_12_20_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_12_20_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_12_20_7  (
            .in0(N__33049),
            .in1(N__33519),
            .in2(_gnd_net_),
            .in3(N__30659),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48341),
            .ce(),
            .sr(N__47838));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_29_LC_12_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_29_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_29_LC_12_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_29_LC_12_21_3  (
            .in0(N__30623),
            .in1(N__30647),
            .in2(_gnd_net_),
            .in3(N__33318),
            .lcout(\delay_measurement_inst.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_12_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_12_21_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__30598),
            .in2(_gnd_net_),
            .in3(N__30622),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_12_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_12_22_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_12_22_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_12_22_4  (
            .in0(N__30605),
            .in1(N__33473),
            .in2(_gnd_net_),
            .in3(N__33127),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48335),
            .ce(),
            .sr(N__47854));
    defparam SB_DFF_inst_DELAY_HC1_LC_13_2_3.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_2_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_13_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30587),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48466),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_13_2_7.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_13_2_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_13_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_13_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30575),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48466),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_13_3_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_13_3_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_13_3_2  (
            .in0(N__30821),
            .in1(N__30791),
            .in2(N__30809),
            .in3(N__30800),
            .lcout(\phase_controller_inst1.stoper_tr.N_248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_13_3_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_13_3_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_13_3_4  (
            .in0(N__38241),
            .in1(N__38686),
            .in2(N__38471),
            .in3(N__34864),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_13_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_13_3_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_13_3_5  (
            .in0(_gnd_net_),
            .in1(N__35064),
            .in2(_gnd_net_),
            .in3(N__35037),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_3_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_3_6 .LUT_INIT=16'b1101110011011101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_3_6  (
            .in0(N__38453),
            .in1(N__38545),
            .in2(N__30794),
            .in3(N__38687),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_4_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_4_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_4_0 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_4_0  (
            .in0(N__40834),
            .in1(N__40935),
            .in2(N__41428),
            .in3(N__37273),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48447),
            .ce(N__30871),
            .sr(N__47747));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_13_4_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_13_4_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_13_4_3  (
            .in0(N__34971),
            .in1(N__35169),
            .in2(_gnd_net_),
            .in3(N__35133),
            .lcout(\phase_controller_inst1.stoper_tr.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_13_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_13_5_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_13_5_1  (
            .in0(N__39205),
            .in1(N__39327),
            .in2(_gnd_net_),
            .in3(N__34998),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_13_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_13_5_2 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(N__38462),
            .in2(N__30782),
            .in3(N__35038),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_5_3 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_13_5_3  (
            .in0(_gnd_net_),
            .in1(N__34860),
            .in2(N__30779),
            .in3(N__38046),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48439),
            .ce(N__42701),
            .sr(N__47753));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_13_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_13_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_13_5_7 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_13_5_7  (
            .in0(N__38285),
            .in1(N__38045),
            .in2(N__35113),
            .in3(N__34938),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48439),
            .ce(N__42701),
            .sr(N__47753));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_13_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_13_6_0 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_13_6_0  (
            .in0(N__40928),
            .in1(N__40983),
            .in2(N__30889),
            .in3(N__41121),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_13_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_13_6_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_13_6_1 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_13_6_1  (
            .in0(N__30933),
            .in1(N__40700),
            .in2(N__39259),
            .in3(N__40775),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48430),
            .ce(N__30872),
            .sr(N__47758));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_13_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_13_6_2 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_13_6_2  (
            .in0(N__40696),
            .in1(N__39252),
            .in2(N__40727),
            .in3(N__30935),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48430),
            .ce(N__30872),
            .sr(N__47758));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_13_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_13_6_4 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_13_6_4  (
            .in0(N__40748),
            .in1(N__39251),
            .in2(N__40703),
            .in3(N__30934),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48430),
            .ce(N__30872),
            .sr(N__47758));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_13_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_13_6_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_13_6_6  (
            .in0(N__38117),
            .in1(N__38129),
            .in2(N__41456),
            .in3(N__30839),
            .lcout(\delay_measurement_inst.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_7_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_7_1  (
            .in0(N__41112),
            .in1(N__40691),
            .in2(N__45650),
            .in3(N__40771),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_7_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_7_2  (
            .in0(N__40976),
            .in1(N__45594),
            .in2(N__30842),
            .in3(N__40793),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_13_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_13_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__41471),
            .in2(_gnd_net_),
            .in3(N__41486),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_13_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_13_7_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_13_7_5  (
            .in0(N__30833),
            .in1(N__40847),
            .in2(N__41405),
            .in3(N__30827),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_13_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_13_7_6 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_13_7_6  (
            .in0(N__30927),
            .in1(N__40833),
            .in2(N__30902),
            .in3(N__30899),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_13_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_13_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_13_7_7  (
            .in0(N__38706),
            .in1(N__35085),
            .in2(N__38583),
            .in3(N__38359),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_13_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_13_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__38611),
            .in2(_gnd_net_),
            .in3(N__35092),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48410),
            .ce(N__42700),
            .sr(N__47771));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_13_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_13_8_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_13_8_4  (
            .in0(N__38612),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38713),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48410),
            .ce(N__42700),
            .sr(N__47771));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_13_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_13_8_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_13_8_6  (
            .in0(N__38551),
            .in1(N__38472),
            .in2(_gnd_net_),
            .in3(N__38688),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_13_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_13_8_7 .LUT_INIT=16'b1010111010101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_13_8_7  (
            .in0(N__35065),
            .in1(N__38497),
            .in2(N__30893),
            .in3(N__35033),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48410),
            .ce(N__42700),
            .sr(N__47771));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_9_0 .LUT_INIT=16'b0000010110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_9_0  (
            .in0(N__36376),
            .in1(N__36608),
            .in2(N__36872),
            .in3(N__36332),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48403),
            .ce(N__35920),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_13_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_13_9_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_0_LC_13_9_1  (
            .in0(N__37440),
            .in1(N__37730),
            .in2(N__37665),
            .in3(N__38176),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48403),
            .ce(N__35920),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_13_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_13_9_2 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_1_LC_13_9_2  (
            .in0(N__38177),
            .in1(N__37618),
            .in2(N__37784),
            .in3(N__37441),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48403),
            .ce(N__35920),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_13_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_13_10_0 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_13_10_0  (
            .in0(N__31400),
            .in1(N__31293),
            .in2(N__31268),
            .in3(N__31226),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_13_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_13_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_13_10_1  (
            .in0(N__31204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31395),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_13_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_13_10_2 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_13_10_2  (
            .in0(N__31401),
            .in1(N__31190),
            .in2(N__31145),
            .in3(N__31142),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_10_3  (
            .in0(N__31116),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31396),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_13_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_13_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_13_10_4  (
            .in0(N__31398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31086),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_6  (
            .in0(N__31397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31062),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_13_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_13_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_13_10_7  (
            .in0(N__31035),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31399),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_13_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_13_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_13_11_0  (
            .in0(N__31640),
            .in1(N__31013),
            .in2(N__31001),
            .in3(N__30986),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_13_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_13_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31682),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_13_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_13_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31917),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEC8M_18_LC_13_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEC8M_18_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEC8M_18_LC_13_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEC8M_18_LC_13_11_3  (
            .in0(N__31847),
            .in1(N__31784),
            .in2(N__31744),
            .in3(N__31683),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_11_4  (
            .in0(N__31630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31392),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_13_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_13_11_5 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_13_11_5  (
            .in0(N__31394),
            .in1(N__31615),
            .in2(N__31571),
            .in3(N__31568),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_13_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_13_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_13_11_6  (
            .in0(N__31539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31391),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_11_7  (
            .in0(N__31393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31294),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__32537),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__31274),
            .in2(N__32831),
            .in3(N__35679),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__32090),
            .in2(N__33818),
            .in3(N__32101),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__32069),
            .in2(N__32744),
            .in3(N__32080),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_12_4  (
            .in0(N__32062),
            .in1(N__32051),
            .in2(N__32381),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_12_5  (
            .in0(N__32044),
            .in1(N__32033),
            .in2(N__32327),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__32000),
            .in2(N__32027),
            .in3(N__32011),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_12_7  (
            .in0(N__31993),
            .in1(N__31982),
            .in2(N__32693),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__31961),
            .in2(N__32621),
            .in3(N__31972),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__31925),
            .in2(N__31955),
            .in3(N__31936),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__32180),
            .in2(N__32594),
            .in3(N__35644),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__32174),
            .in2(N__32609),
            .in3(N__35719),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_13_4  (
            .in0(N__32237),
            .in1(N__32168),
            .in2(N__32312),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__32162),
            .in2(N__34442),
            .in3(N__32216),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__32141),
            .in2(N__32156),
            .in3(N__32195),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__32135),
            .in2(N__34379),
            .in3(N__32522),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__32129),
            .in2(N__32888),
            .in3(N__32500),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__32111),
            .in2(N__32123),
            .in3(N__32482),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__32282),
            .in2(N__32297),
            .in3(N__32464),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__32276),
            .in2(N__36089),
            .in3(N__32446),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32270),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36704),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35936),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_13_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_13_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__35826),
            .in2(_gnd_net_),
            .in3(N__35781),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_15_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_15_0  (
            .in0(N__36472),
            .in1(N__36319),
            .in2(N__36601),
            .in3(N__32243),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_15_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_15_1  (
            .in0(N__36315),
            .in1(N__36551),
            .in2(N__36478),
            .in3(N__32222),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_15_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_15_2  (
            .in0(N__36473),
            .in1(N__36320),
            .in2(N__36602),
            .in3(N__32201),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_15_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_15_3  (
            .in0(N__36316),
            .in1(N__36552),
            .in2(N__36479),
            .in3(N__32528),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_15_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_15_4  (
            .in0(N__36474),
            .in1(N__36321),
            .in2(N__36603),
            .in3(N__32507),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_15_5 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_15_5  (
            .in0(N__36317),
            .in1(N__32489),
            .in2(N__36481),
            .in3(N__36566),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_15_6 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_15_6  (
            .in0(N__36475),
            .in1(N__32471),
            .in2(N__36604),
            .in3(N__36322),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_15_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_15_7  (
            .in0(N__36318),
            .in1(N__36553),
            .in2(N__36480),
            .in3(N__32453),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48373),
            .ce(),
            .sr(N__47801));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_13_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_13_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_13_16_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_13_16_0  (
            .in0(N__34294),
            .in1(N__32435),
            .in2(N__33959),
            .in3(N__34166),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_13_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_13_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_13_16_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_13_16_1  (
            .in0(N__34167),
            .in1(N__32365),
            .in2(N__34337),
            .in3(N__33910),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_13_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_13_16_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_13_16_2  (
            .in0(N__34293),
            .in1(N__33755),
            .in2(N__33958),
            .in3(N__34165),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_13_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_13_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_13_16_3 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_13_16_3  (
            .in0(N__32934),
            .in1(N__33908),
            .in2(_gnd_net_),
            .in3(N__34296),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_13_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_13_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_13_16_4 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_13_16_4  (
            .in0(N__33907),
            .in1(N__32876),
            .in2(_gnd_net_),
            .in3(N__32816),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5  (
            .in0(N__32817),
            .in1(N__33909),
            .in2(_gnd_net_),
            .in3(N__32794),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_13_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_13_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_13_16_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_13_16_6  (
            .in0(N__34295),
            .in1(N__32732),
            .in2(N__33960),
            .in3(N__34168),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_13_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_13_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_13_16_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_13_16_7  (
            .in0(N__34169),
            .in1(N__32678),
            .in2(N__34338),
            .in3(N__33911),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48368),
            .ce(N__36075),
            .sr(N__47805));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_13_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_13_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_13_17_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_13_17_0  (
            .in0(N__34172),
            .in1(N__33704),
            .in2(N__33962),
            .in3(N__34268),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48364),
            .ce(N__36077),
            .sr(N__47810));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_17_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_13_17_1  (
            .in0(N__34265),
            .in1(N__33927),
            .in2(N__33593),
            .in3(N__34171),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48364),
            .ce(N__36077),
            .sr(N__47810));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_17_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_17_2  (
            .in0(N__36147),
            .in1(N__32579),
            .in2(N__36207),
            .in3(N__36130),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_13_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_13_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_13_17_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_0_LC_13_17_3  (
            .in0(N__34264),
            .in1(N__34170),
            .in2(N__32573),
            .in3(N__32570),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48364),
            .ce(N__36077),
            .sr(N__47810));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_13_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_13_17_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_13_17_5  (
            .in0(N__34266),
            .in1(N__33928),
            .in2(N__34508),
            .in3(N__34173),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48364),
            .ce(N__36077),
            .sr(N__47810));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_13_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_13_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_13_17_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_13_17_6  (
            .in0(N__34174),
            .in1(N__34430),
            .in2(N__33963),
            .in3(N__34269),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48364),
            .ce(N__36077),
            .sr(N__47810));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_13_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_13_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_13_17_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_13_17_7  (
            .in0(N__34267),
            .in1(N__34175),
            .in2(N__34054),
            .in3(N__33935),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48364),
            .ce(N__36077),
            .sr(N__47810));
    defparam \phase_controller_inst1.state_3_LC_13_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_18_7 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_18_7  (
            .in0(N__33803),
            .in1(N__43856),
            .in2(N__34611),
            .in3(N__33773),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48358),
            .ce(),
            .sr(N__47815));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_20_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_20_2  (
            .in0(N__33751),
            .in1(N__33702),
            .in2(N__33642),
            .in3(N__33574),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_21_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_21_3 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_13_21_3  (
            .in0(N__33515),
            .in1(N__33319),
            .in2(N__32967),
            .in3(N__33128),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48343),
            .ce(),
            .sr(N__47839));
    defparam \current_shift_inst.timer_s1.running_LC_13_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_25_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_25_1  (
            .in0(N__36983),
            .in1(N__37004),
            .in2(_gnd_net_),
            .in3(N__34547),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48332),
            .ce(),
            .sr(N__47867));
    defparam \phase_controller_inst1.S1_LC_13_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34610),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48332),
            .ce(),
            .sr(N__47867));
    defparam \current_shift_inst.start_timer_s1_LC_13_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_25_3 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_25_3  (
            .in0(N__34608),
            .in1(N__34560),
            .in2(_gnd_net_),
            .in3(N__34545),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48332),
            .ce(),
            .sr(N__47867));
    defparam \current_shift_inst.stop_timer_s1_LC_13_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_25_6 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_25_6  (
            .in0(N__34546),
            .in1(N__34609),
            .in2(N__34567),
            .in3(N__36982),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48332),
            .ce(),
            .sr(N__47867));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_26_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_26_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_26_7  (
            .in0(N__37001),
            .in1(N__36980),
            .in2(_gnd_net_),
            .in3(N__34544),
            .lcout(\current_shift_inst.timer_s1.N_181_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_27_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_27_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43380),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48329),
            .ce(),
            .sr(N__47876));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_2_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_2_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_2_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_2_1  (
            .in0(N__37786),
            .in1(N__37677),
            .in2(N__37529),
            .in3(N__37151),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48471),
            .ce(),
            .sr(N__47735));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_14_2_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_14_2_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(N__37518),
            .in2(_gnd_net_),
            .in3(N__37785),
            .lcout(\phase_controller_inst2.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst2.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_2_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_2_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_2_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34511),
            .in3(N__38181),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_3_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_3_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_3_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_3_0  (
            .in0(N__37792),
            .in1(N__37683),
            .in2(N__37355),
            .in3(N__37491),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48467),
            .ce(),
            .sr(N__47738));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_3_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_3_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_3_2 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_3_2  (
            .in0(N__37791),
            .in1(N__37682),
            .in2(N__37016),
            .in3(N__37490),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48467),
            .ce(),
            .sr(N__47738));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_3_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_3_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_3_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_3_6  (
            .in0(N__37790),
            .in1(N__37681),
            .in2(N__37097),
            .in3(N__37489),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48467),
            .ce(),
            .sr(N__47738));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_3_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_3_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_3_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_3_7  (
            .in0(N__37488),
            .in1(N__37793),
            .in2(N__37685),
            .in3(N__36935),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48467),
            .ce(),
            .sr(N__47738));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_4_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_4_0  (
            .in0(N__37788),
            .in1(N__37527),
            .in2(N__37672),
            .in3(N__37301),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__47740));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_4_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_4_1  (
            .in0(N__37524),
            .in1(N__37630),
            .in2(N__37812),
            .in3(N__37067),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__47740));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_4_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_4_4  (
            .in0(N__37789),
            .in1(N__37528),
            .in2(N__37673),
            .in3(N__37127),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__47740));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_4_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_4_6  (
            .in0(N__37787),
            .in1(N__37526),
            .in2(N__37671),
            .in3(N__37043),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__47740));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_4_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_4_7  (
            .in0(N__37525),
            .in1(N__37631),
            .in2(N__37813),
            .in3(N__37325),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__47740));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38749),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(N__42705),
            .sr(N__47748));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_14_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_14_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_14_5_2 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_14_5_2  (
            .in0(N__38275),
            .in1(N__38101),
            .in2(_gnd_net_),
            .in3(N__35008),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(N__42705),
            .sr(N__47748));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_14_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_14_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_14_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_14_5_3  (
            .in0(N__38100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39206),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(N__42705),
            .sr(N__47748));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_14_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_14_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_14_5_6 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_14_5_6  (
            .in0(N__38276),
            .in1(N__34978),
            .in2(N__38105),
            .in3(N__34939),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(N__42705),
            .sr(N__47748));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_14_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_14_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_14_5_7 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_14_5_7  (
            .in0(N__38099),
            .in1(N__38274),
            .in2(N__35170),
            .in3(N__35140),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(N__42705),
            .sr(N__47748));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_14_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_14_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__34730),
            .in2(N__34724),
            .in3(N__37830),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_14_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_14_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__34703),
            .in2(N__34715),
            .in3(N__37957),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_14_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_14_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__34685),
            .in2(N__34697),
            .in3(N__37930),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_14_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_14_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__34679),
            .in2(N__38222),
            .in3(N__36950),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_14_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_14_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__34673),
            .in2(N__34667),
            .in3(N__37906),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_14_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_14_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__34643),
            .in2(N__34658),
            .in3(N__37876),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_14_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_14_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_14_6_6  (
            .in0(N__37180),
            .in1(N__34622),
            .in2(N__34637),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_14_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_14_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__34829),
            .in2(N__34841),
            .in3(N__37169),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_14_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_14_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__34811),
            .in2(N__34823),
            .in3(N__37142),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_14_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_14_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_14_7_1  (
            .in0(N__37852),
            .in1(N__34805),
            .in2(N__38348),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_14_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_14_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__34790),
            .in2(N__34799),
            .in3(N__37381),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_14_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_14_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__34769),
            .in2(N__34784),
            .in3(N__37112),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_14_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_14_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__34763),
            .in2(N__38339),
            .in3(N__37082),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_14_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_14_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__34757),
            .in2(N__38327),
            .in3(N__37058),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_14_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_14_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__34736),
            .in2(N__34751),
            .in3(N__37034),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_14_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_14_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__34922),
            .in2(N__42728),
            .in3(N__37370),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_14_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_14_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__34916),
            .in2(N__34883),
            .in3(N__37343),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_14_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_14_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__34910),
            .in2(N__34874),
            .in3(N__37316),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_14_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_14_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__34892),
            .in2(N__34904),
            .in3(N__37214),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34886),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39127),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48421),
            .ce(N__42709),
            .sr(N__47767));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39079),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48421),
            .ce(N__42709),
            .sr(N__47767));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_14_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_14_9_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_14_9_2  (
            .in0(N__38312),
            .in1(N__38096),
            .in2(_gnd_net_),
            .in3(N__38249),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48411),
            .ce(N__39037),
            .sr(N__47772));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_14_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_14_9_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_14_9_3  (
            .in0(N__38094),
            .in1(N__34865),
            .in2(_gnd_net_),
            .in3(N__38313),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48411),
            .ce(N__39037),
            .sr(N__47772));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_14_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_14_9_4 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_14_9_4  (
            .in0(N__38311),
            .in1(N__38095),
            .in2(N__35177),
            .in3(N__35144),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48411),
            .ce(N__39037),
            .sr(N__47772));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_14_9_6 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_14_9_6  (
            .in0(N__38314),
            .in1(N__38097),
            .in2(N__35120),
            .in3(N__34951),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48411),
            .ce(N__39037),
            .sr(N__47772));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_14_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_14_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_14_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__38093),
            .in2(_gnd_net_),
            .in3(N__39331),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_14_10_1  (
            .in0(N__38626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38375),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_14_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__38627),
            .in2(_gnd_net_),
            .in3(N__35096),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_14_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_14_10_3 .LUT_INIT=16'b1010111010101111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_14_10_3  (
            .in0(N__35069),
            .in1(N__38499),
            .in2(N__38641),
            .in3(N__35039),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_14_10_4 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_14_10_4  (
            .in0(N__35009),
            .in1(N__38092),
            .in2(_gnd_net_),
            .in3(N__38307),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_14_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_14_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_14_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42764),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_14_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_14_10_7 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_14_10_7  (
            .in0(N__38091),
            .in1(N__34982),
            .in2(N__38315),
            .in3(N__34952),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(N__39036),
            .sr(N__47777));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_11_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_11_0  (
            .in0(N__43562),
            .in1(N__43818),
            .in2(N__43717),
            .in3(N__41975),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_11_1  (
            .in0(N__43914),
            .in1(N__41329),
            .in2(_gnd_net_),
            .in3(N__43882),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_2  (
            .in0(N__43565),
            .in1(N__43696),
            .in2(N__35180),
            .in3(N__43821),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_11_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_11_3  (
            .in0(N__43815),
            .in1(N__43687),
            .in2(N__43575),
            .in3(N__41942),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_11_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_11_4  (
            .in0(N__43563),
            .in1(N__43819),
            .in2(N__43718),
            .in3(N__41909),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_11_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_11_5  (
            .in0(N__43816),
            .in1(N__43691),
            .in2(N__43576),
            .in3(N__41876),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_11_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_11_6  (
            .in0(N__43564),
            .in1(N__43820),
            .in2(N__43719),
            .in3(N__41843),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_11_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_11_7  (
            .in0(N__43817),
            .in1(N__43695),
            .in2(N__43577),
            .in3(N__41810),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(N__47779));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_12_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_12_0  (
            .in0(N__43776),
            .in1(N__43630),
            .in2(N__43554),
            .in3(N__41600),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48393),
            .ce(),
            .sr(N__47786));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_12_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_12_1  (
            .in0(N__43517),
            .in1(N__43778),
            .in2(N__43660),
            .in3(N__41561),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48393),
            .ce(),
            .sr(N__47786));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_12_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_12_2  (
            .in0(N__43777),
            .in1(N__43634),
            .in2(N__43555),
            .in3(N__41531),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48393),
            .ce(),
            .sr(N__47786));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_12_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_12_3  (
            .in0(N__43629),
            .in1(N__43506),
            .in2(_gnd_net_),
            .in3(N__43775),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_14_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_14_12_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_14_12_4  (
            .in0(N__36916),
            .in1(N__35683),
            .in2(_gnd_net_),
            .in3(N__36861),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_12_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_12_5  (
            .in0(N__36579),
            .in1(N__36446),
            .in2(N__35693),
            .in3(N__36288),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48393),
            .ce(),
            .sr(N__47786));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_7  (
            .in0(N__36463),
            .in1(N__36287),
            .in2(N__36609),
            .in3(N__35663),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48393),
            .ce(),
            .sr(N__47786));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_14_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_14_13_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_14_13_0  (
            .in0(N__35214),
            .in1(N__35355),
            .in2(N__35585),
            .in3(N__35632),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_14_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_14_13_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_14_13_1  (
            .in0(N__35633),
            .in1(N__35574),
            .in2(N__35375),
            .in3(N__35215),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_13_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_13_3  (
            .in0(N__43518),
            .in1(N__43804),
            .in2(N__43724),
            .in3(N__43880),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_13_4 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_13_4  (
            .in0(N__43881),
            .in1(N__43716),
            .in2(N__43823),
            .in3(N__43519),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__43915),
            .in2(_gnd_net_),
            .in3(N__43878),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_13_6  (
            .in0(N__43879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43916),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_14_13_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_0_LC_14_13_7  (
            .in0(N__36459),
            .in1(N__36289),
            .in2(N__36605),
            .in3(N__36860),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_14_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_14_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__35745),
            .in2(_gnd_net_),
            .in3(N__36807),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_hc_RNO_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_14_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_14_14_1 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_14_14_1  (
            .in0(N__35843),
            .in1(N__36550),
            .in2(N__35834),
            .in3(N__45481),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48385),
            .ce(),
            .sr(N__47793));
    defparam \phase_controller_inst2.state_2_LC_14_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_14_14_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_2_LC_14_14_3  (
            .in0(N__36808),
            .in1(N__35827),
            .in2(N__35752),
            .in3(N__35785),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48385),
            .ce(),
            .sr(N__47793));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_14_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_14_4  (
            .in0(N__36549),
            .in1(N__36254),
            .in2(N__36482),
            .in3(N__35732),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48385),
            .ce(),
            .sr(N__47793));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_14_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_14_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__36427),
            .in2(_gnd_net_),
            .in3(N__36253),
            .lcout(\phase_controller_inst2.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_inst2.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_14_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35708),
            .in3(N__36849),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_14_15_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_14_15_0  (
            .in0(N__36212),
            .in1(N__36155),
            .in2(_gnd_net_),
            .in3(N__36131),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48379),
            .ce(N__36062),
            .sr(N__47797));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_15_2  (
            .in0(N__36785),
            .in1(_gnd_net_),
            .in2(N__45966),
            .in3(N__45434),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_15_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__45907),
            .in2(N__36029),
            .in3(N__42064),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_14_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_14_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__36903),
            .in2(_gnd_net_),
            .in3(N__36850),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_0_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_14_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__39167),
            .in2(N__39161),
            .in3(N__39160),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_14_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__39146),
            .in2(_gnd_net_),
            .in3(N__35975),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_14_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__39140),
            .in2(_gnd_net_),
            .in3(N__35954),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_14_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__39407),
            .in2(_gnd_net_),
            .in3(N__35939),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_14_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__39401),
            .in2(_gnd_net_),
            .in3(N__36743),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_14_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__39395),
            .in2(_gnd_net_),
            .in3(N__36728),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_14_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__39389),
            .in2(_gnd_net_),
            .in3(N__36707),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_14_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__39359),
            .in2(_gnd_net_),
            .in3(N__36692),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__48374),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__36758),
            .in2(_gnd_net_),
            .in3(N__36671),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__48369),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_14_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__39353),
            .in2(_gnd_net_),
            .in3(N__36659),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__48369),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_14_17_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_10_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39344),
            .in3(N__36656),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__48369),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_14_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_11_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_14_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.control_input_11_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__39662),
            .in2(_gnd_net_),
            .in3(N__36653),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48369),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_17_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_17_4  (
            .in0(N__36607),
            .in1(N__36476),
            .in2(_gnd_net_),
            .in3(N__36296),
            .lcout(\phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_17_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_17_5  (
            .in0(N__49581),
            .in1(N__36752),
            .in2(_gnd_net_),
            .in3(N__48512),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_17_6  (
            .in0(N__36776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_17_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_17_7  (
            .in0(N__46462),
            .in1(N__42224),
            .in2(_gnd_net_),
            .in3(N__39521),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_0  (
            .in0(N__49566),
            .in1(N__47137),
            .in2(N__49280),
            .in3(N__47102),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48722),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48365),
            .ce(N__47988),
            .sr(N__47811));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_18_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_18_3  (
            .in0(N__46961),
            .in1(N__49565),
            .in2(N__49281),
            .in3(N__46193),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_18_4 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_18_4  (
            .in0(N__46192),
            .in1(N__49110),
            .in2(N__49645),
            .in3(N__46962),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45325),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_18_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__49561),
            .in2(N__36746),
            .in3(N__48508),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_0  (
            .in0(N__49580),
            .in1(N__46545),
            .in2(N__49394),
            .in3(N__46505),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_19_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_19_1  (
            .in0(N__49588),
            .in1(N__49309),
            .in2(N__42500),
            .in3(N__45020),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2  (
            .in0(N__49579),
            .in1(N__46926),
            .in2(N__49393),
            .in3(N__46886),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_19_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_19_3  (
            .in0(N__49590),
            .in1(N__49311),
            .in2(N__46783),
            .in3(N__46736),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_19_4  (
            .in0(N__49578),
            .in1(N__46854),
            .in2(N__49395),
            .in3(N__46814),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_19_5 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_19_5  (
            .in0(N__49589),
            .in1(N__47066),
            .in2(N__44957),
            .in3(N__49310),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_19_6  (
            .in0(N__49577),
            .in1(N__44161),
            .in2(N__49396),
            .in3(N__44465),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_19_7 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_19_7  (
            .in0(N__49587),
            .in1(N__44416),
            .in2(N__44675),
            .in3(N__49308),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_14_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_14_21_0 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_14_21_0  (
            .in0(N__36806),
            .in1(N__36917),
            .in2(N__36887),
            .in3(N__36868),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48347),
            .ce(),
            .sr(N__47830));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48705),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48338),
            .ce(N__47954),
            .sr(N__47848));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_25_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__37002),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_14_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_14_25_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_14_25_1  (
            .in0(N__37003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36981),
            .lcout(\current_shift_inst.timer_s1.N_180_i_g ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_2_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_2_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_2_0  (
            .in0(_gnd_net_),
            .in1(N__36962),
            .in2(N__37838),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_2_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_15_2_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_15_2_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_15_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_15_2_1  (
            .in0(_gnd_net_),
            .in1(N__37961),
            .in2(_gnd_net_),
            .in3(N__36956),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_15_2_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_15_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_15_2_2  (
            .in0(_gnd_net_),
            .in1(N__38141),
            .in2(N__37937),
            .in3(N__36953),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_15_2_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_15_2_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_15_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_15_2_3  (
            .in0(_gnd_net_),
            .in1(N__36949),
            .in2(_gnd_net_),
            .in3(N__36929),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_15_2_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_15_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(N__37910),
            .in2(_gnd_net_),
            .in3(N__36926),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_15_2_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_15_2_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_15_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_15_2_5  (
            .in0(_gnd_net_),
            .in1(N__37883),
            .in2(_gnd_net_),
            .in3(N__36923),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_15_2_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_15_2_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_15_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_15_2_6  (
            .in0(_gnd_net_),
            .in1(N__37184),
            .in2(_gnd_net_),
            .in3(N__36920),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_15_2_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_15_2_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_15_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_15_2_7  (
            .in0(_gnd_net_),
            .in1(N__37165),
            .in2(_gnd_net_),
            .in3(N__37145),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_15_3_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_15_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(N__37141),
            .in2(_gnd_net_),
            .in3(N__37121),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_15_3_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_15_3_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_15_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_15_3_1  (
            .in0(_gnd_net_),
            .in1(N__37856),
            .in2(_gnd_net_),
            .in3(N__37118),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_15_3_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_15_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_15_3_2  (
            .in0(_gnd_net_),
            .in1(N__37385),
            .in2(_gnd_net_),
            .in3(N__37115),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_15_3_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_15_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_15_3_3  (
            .in0(_gnd_net_),
            .in1(N__37111),
            .in2(_gnd_net_),
            .in3(N__37085),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_15_3_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_15_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_15_3_4  (
            .in0(_gnd_net_),
            .in1(N__37081),
            .in2(_gnd_net_),
            .in3(N__37061),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_15_3_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_15_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(N__37057),
            .in2(_gnd_net_),
            .in3(N__37037),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_15_3_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_15_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(N__37030),
            .in2(_gnd_net_),
            .in3(N__37007),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_15_3_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_15_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_15_3_7  (
            .in0(_gnd_net_),
            .in1(N__37369),
            .in2(_gnd_net_),
            .in3(N__37346),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_15_4_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_15_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__37339),
            .in2(_gnd_net_),
            .in3(N__37319),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_15_4_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_15_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__37315),
            .in2(_gnd_net_),
            .in3(N__37295),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_15_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_15_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__37210),
            .in2(_gnd_net_),
            .in3(N__37292),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_4_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_4_4 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_4_4  (
            .in0(N__40829),
            .in1(N__37289),
            .in2(N__41417),
            .in3(N__37274),
            .lcout(\delay_measurement_inst.N_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_15_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_15_4_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_15_4_6  (
            .in0(N__37622),
            .in1(N__37523),
            .in2(_gnd_net_),
            .in3(N__37814),
            .lcout(\phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_5_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_5_0  (
            .in0(N__37512),
            .in1(N__37803),
            .in2(N__37674),
            .in3(N__37220),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_5_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_5_1  (
            .in0(N__37802),
            .in1(N__37652),
            .in2(N__37196),
            .in3(N__37517),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_15_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_15_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_15_5_2 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_15_5_2  (
            .in0(N__37989),
            .in1(N__38208),
            .in2(N__38009),
            .in3(N__38183),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_5_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_5_3  (
            .in0(N__37800),
            .in1(N__37650),
            .in2(N__37973),
            .in3(N__37515),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_5_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_5_4  (
            .in0(N__37513),
            .in1(N__37804),
            .in2(N__37675),
            .in3(N__37946),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_5_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_5_6  (
            .in0(N__37514),
            .in1(N__37805),
            .in2(N__37676),
            .in3(N__37919),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_5_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_5_7  (
            .in0(N__37801),
            .in1(N__37651),
            .in2(N__37895),
            .in3(N__37516),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__47741));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_6_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_6_0  (
            .in0(N__37492),
            .in1(N__37810),
            .in2(N__37684),
            .in3(N__37865),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(),
            .sr(N__47749));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_15_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_15_6_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_15_6_1  (
            .in0(N__38210),
            .in1(N__37834),
            .in2(_gnd_net_),
            .in3(N__38182),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_15_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_15_6_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_15_6_2  (
            .in0(N__37666),
            .in1(N__37493),
            .in2(N__37841),
            .in3(N__37811),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(),
            .sr(N__47749));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_6_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_6_3  (
            .in0(N__37809),
            .in1(N__37667),
            .in2(N__37522),
            .in3(N__37394),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(),
            .sr(N__47749));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_7_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_15_7_2  (
            .in0(N__38371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38642),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48440),
            .ce(N__42687),
            .sr(N__47754));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_15_7_3  (
            .in0(N__38643),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38590),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48440),
            .ce(N__42687),
            .sr(N__47754));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_15_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_15_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_15_7_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_15_7_5  (
            .in0(N__38550),
            .in1(N__38498),
            .in2(_gnd_net_),
            .in3(N__38692),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48440),
            .ce(N__42687),
            .sr(N__47754));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_15_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_15_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_15_7_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_15_7_6  (
            .in0(N__38297),
            .in1(N__38098),
            .in2(_gnd_net_),
            .in3(N__38248),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48440),
            .ce(N__42687),
            .sr(N__47754));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_15_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__38209),
            .in2(_gnd_net_),
            .in3(N__38172),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_15_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_15_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_15_8_1  (
            .in0(N__41510),
            .in1(N__41519),
            .in2(N__41501),
            .in3(N__41162),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_15_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_15_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_15_8_3  (
            .in0(N__41183),
            .in1(N__41192),
            .in2(N__41174),
            .in3(N__41201),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42589),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__38068),
            .in2(_gnd_net_),
            .in3(N__39204),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(N__39038),
            .sr(N__47768));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38753),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(N__39038),
            .sr(N__47768));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__38644),
            .in2(_gnd_net_),
            .in3(N__38717),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(N__39038),
            .sr(N__47768));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_9_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_15_9_4  (
            .in0(N__38693),
            .in1(N__38557),
            .in2(_gnd_net_),
            .in3(N__38501),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(N__39038),
            .sr(N__47768));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__38645),
            .in2(_gnd_net_),
            .in3(N__38591),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(N__39038),
            .sr(N__47768));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__38558),
            .in2(_gnd_net_),
            .in3(N__38500),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(N__39038),
            .sr(N__47768));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__38411),
            .in2(N__38420),
            .in3(N__41319),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__38396),
            .in2(N__38405),
            .in3(N__41305),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__38381),
            .in2(N__38390),
            .in3(N__41743),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__38870),
            .in2(N__38882),
            .in3(N__41713),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__38852),
            .in2(N__38864),
            .in3(N__41683),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__38837),
            .in2(N__38846),
            .in3(N__41650),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__38822),
            .in2(N__38831),
            .in3(N__41617),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__38804),
            .in2(N__38816),
            .in3(N__41584),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__38789),
            .in2(N__38798),
            .in3(N__41542),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_11_1  (
            .in0(N__41986),
            .in1(N__38774),
            .in2(N__38783),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__38759),
            .in2(N__38768),
            .in3(N__41953),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__38993),
            .in2(N__39005),
            .in3(N__41920),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__38975),
            .in2(N__38987),
            .in3(N__41887),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__38954),
            .in2(N__38969),
            .in3(N__41854),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__38936),
            .in2(N__38948),
            .in3(N__41821),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_11_7  (
            .in0(N__43931),
            .in1(N__38921),
            .in2(N__38930),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__38915),
            .in2(N__39092),
            .in3(N__41791),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__38909),
            .in2(N__39047),
            .in3(N__42109),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__38888),
            .in2(N__38903),
            .in3(N__42088),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39134),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39131),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48398),
            .ce(N__39026),
            .sr(N__47780));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39083),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48398),
            .ce(N__39026),
            .sr(N__47780));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_13_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_13_0  (
            .in0(N__43513),
            .in1(N__43797),
            .in2(N__43720),
            .in3(N__41780),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_13_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_13_1  (
            .in0(N__43794),
            .in1(N__43700),
            .in2(N__43556),
            .in3(N__42098),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_13_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_13_2  (
            .in0(N__43514),
            .in1(N__43798),
            .in2(N__43721),
            .in3(N__42074),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_13_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_13_3  (
            .in0(N__43795),
            .in1(N__43704),
            .in2(N__43557),
            .in3(N__41771),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_13_4 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_13_4  (
            .in0(N__41726),
            .in1(N__43526),
            .in2(N__43722),
            .in3(N__43800),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_13_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_13_5  (
            .in0(N__43796),
            .in1(N__43708),
            .in2(N__43558),
            .in3(N__41696),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_13_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_13_6  (
            .in0(N__43515),
            .in1(N__43799),
            .in2(N__43723),
            .in3(N__41666),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_13_7 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_13_7  (
            .in0(N__41633),
            .in1(N__43516),
            .in2(N__43822),
            .in3(N__43712),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(N__47787));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46694),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_15_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_15_14_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_15_14_1  (
            .in0(N__45231),
            .in1(N__49741),
            .in2(N__49391),
            .in3(N__44794),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_14_2  (
            .in0(N__49744),
            .in1(N__44412),
            .in2(N__49388),
            .in3(N__44671),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_14_3  (
            .in0(N__48686),
            .in1(N__42492),
            .in2(_gnd_net_),
            .in3(N__45018),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_15_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_15_14_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_15_14_4  (
            .in0(N__45019),
            .in1(N__49292),
            .in2(N__42499),
            .in3(N__49749),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_14_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_14_5  (
            .in0(N__49750),
            .in1(N__47069),
            .in2(N__49390),
            .in3(N__44956),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_6  (
            .in0(N__49743),
            .in1(N__44536),
            .in2(N__49389),
            .in3(N__44627),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_14_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_14_7  (
            .in0(N__45232),
            .in1(N__49742),
            .in2(N__49392),
            .in3(N__44795),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_15_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_15_0  (
            .in0(N__42236),
            .in1(N__39536),
            .in2(_gnd_net_),
            .in3(N__46459),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_15_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_15_2  (
            .in0(N__39509),
            .in1(N__42212),
            .in2(_gnd_net_),
            .in3(N__46460),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_15_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_15_3  (
            .in0(N__46461),
            .in1(N__39497),
            .in2(_gnd_net_),
            .in3(N__42200),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_15_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_15_15_6  (
            .in0(N__39247),
            .in1(N__40637),
            .in2(N__39326),
            .in3(N__39286),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48386),
            .ce(),
            .sr(N__47794));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_15_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_15_15_7  (
            .in0(N__39287),
            .in1(N__39248),
            .in2(N__39189),
            .in3(N__41153),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48386),
            .ce(),
            .sr(N__47794));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_16_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_16_0  (
            .in0(N__39464),
            .in1(N__42167),
            .in2(_gnd_net_),
            .in3(N__46438),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_16_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_16_1  (
            .in0(N__46439),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.N_1318_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_16_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_16_2  (
            .in0(N__39452),
            .in1(N__42158),
            .in2(_gnd_net_),
            .in3(N__46440),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_16_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_16_3  (
            .in0(N__46441),
            .in1(N__39620),
            .in2(_gnd_net_),
            .in3(N__42149),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_16_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_16_4  (
            .in0(N__42140),
            .in1(N__39605),
            .in2(_gnd_net_),
            .in3(N__46442),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_16_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_16_5  (
            .in0(N__46443),
            .in1(N__39581),
            .in2(_gnd_net_),
            .in3(N__42278),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_16_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_16_6  (
            .in0(N__39566),
            .in1(N__42269),
            .in2(_gnd_net_),
            .in3(N__46444),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_16_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_16_7  (
            .in0(N__46445),
            .in1(N__39551),
            .in2(_gnd_net_),
            .in3(N__42260),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__39383),
            .in2(N__42043),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__46403),
            .in2(N__46349),
            .in3(N__45396),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_17_2  (
            .in0(N__45397),
            .in1(N__39377),
            .in2(N__49195),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__48975),
            .in2(N__39371),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__46562),
            .in2(N__49196),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__48979),
            .in2(N__42350),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__39440),
            .in2(N__49197),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__48983),
            .in2(N__42176),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__48984),
            .in2(N__42305),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__48994),
            .in2(N__42359),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__39428),
            .in2(N__49201),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__39422),
            .in2(N__49198),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__42329),
            .in2(N__49202),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__39413),
            .in2(N__49199),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__42395),
            .in2(N__49203),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__39485),
            .in2(N__49200),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__49204),
            .in2(N__42407),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__39479),
            .in2(N__49356),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__49208),
            .in2(N__39473),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__42284),
            .in2(N__49357),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__49212),
            .in2(N__42455),
            .in3(N__39455),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__49802),
            .in2(N__49358),
            .in3(N__39443),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__49216),
            .in2(N__39629),
            .in3(N__39608),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__42386),
            .in2(N__49359),
            .in3(N__39593),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__49220),
            .in2(N__39590),
            .in3(N__39569),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__42365),
            .in2(N__49360),
            .in3(N__39554),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__49224),
            .in2(N__42425),
            .in3(N__39539),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__42461),
            .in2(N__49361),
            .in3(N__39524),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__42371),
            .in2(N__49428),
            .in3(N__39512),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__42446),
            .in2(N__49362),
            .in3(N__39500),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__42439),
            .in2(N__49429),
            .in3(N__39488),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_11_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_11_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_11_LC_15_20_7 .LUT_INIT=16'b1100010100110101;
    LogicCell40 \current_shift_inst.control_input_RNO_0_11_LC_15_20_7  (
            .in0(N__42185),
            .in1(N__49811),
            .in2(N__46466),
            .in3(N__39665),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_21_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__39817),
            .in2(N__48545),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__39796),
            .in2(N__46393),
            .in3(N__39650),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__39818),
            .in2(N__39772),
            .in3(N__39647),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__39797),
            .in2(N__39745),
            .in3(N__39644),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__40039),
            .in2(N__39773),
            .in3(N__39641),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__40015),
            .in2(N__39746),
            .in3(N__39638),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__40040),
            .in2(N__39992),
            .in3(N__39635),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__40016),
            .in2(N__39962),
            .in3(N__39632),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48352),
            .ce(N__48008),
            .sr(N__47822));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__39991),
            .in2(N__39931),
            .in3(N__39692),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__39961),
            .in2(N__39901),
            .in3(N__39689),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__39874),
            .in2(N__39932),
            .in3(N__39686),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__39853),
            .in2(N__39902),
            .in3(N__39683),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__39875),
            .in2(N__40258),
            .in3(N__39680),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__39854),
            .in2(N__40231),
            .in3(N__39677),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__40201),
            .in2(N__40259),
            .in3(N__39674),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__40174),
            .in2(N__40232),
            .in3(N__39671),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48348),
            .ce(N__47995),
            .sr(N__47831));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__40202),
            .in2(N__40144),
            .in3(N__39668),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__40175),
            .in2(N__40114),
            .in3(N__39719),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__40084),
            .in2(N__40145),
            .in3(N__39716),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__40063),
            .in2(N__40115),
            .in3(N__39713),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__40085),
            .in2(N__40609),
            .in3(N__39710),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__40064),
            .in2(N__40579),
            .in3(N__39707),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__40552),
            .in2(N__40610),
            .in3(N__39704),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__40525),
            .in2(N__40580),
            .in3(N__39701),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48344),
            .ce(N__47987),
            .sr(N__47840));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__40553),
            .in2(N__40498),
            .in3(N__39698),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48339),
            .ce(N__47994),
            .sr(N__47849));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__40526),
            .in2(N__40468),
            .in3(N__39695),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48339),
            .ce(N__47994),
            .sr(N__47849));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__40439),
            .in2(N__40499),
            .in3(N__39833),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48339),
            .ce(N__47994),
            .sr(N__47849));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__40295),
            .in2(N__40469),
            .in3(N__39830),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48339),
            .ce(N__47994),
            .sr(N__47849));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39827),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_15_25_0  (
            .in0(N__40380),
            .in1(N__48531),
            .in2(_gnd_net_),
            .in3(N__39824),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_15_25_1  (
            .in0(N__40375),
            .in1(N__46380),
            .in2(_gnd_net_),
            .in3(N__39821),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_15_25_2  (
            .in0(N__40381),
            .in1(N__39816),
            .in2(_gnd_net_),
            .in3(N__39800),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_15_25_3  (
            .in0(N__40376),
            .in1(N__39790),
            .in2(_gnd_net_),
            .in3(N__39776),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_15_25_4  (
            .in0(N__40382),
            .in1(N__39765),
            .in2(_gnd_net_),
            .in3(N__39749),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_15_25_5  (
            .in0(N__40377),
            .in1(N__39738),
            .in2(_gnd_net_),
            .in3(N__39722),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_15_25_6  (
            .in0(N__40379),
            .in1(N__40033),
            .in2(_gnd_net_),
            .in3(N__40019),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_15_25_7  (
            .in0(N__40378),
            .in1(N__40009),
            .in2(_gnd_net_),
            .in3(N__39995),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__48337),
            .ce(N__40277),
            .sr(N__47855));
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_15_26_0  (
            .in0(N__40386),
            .in1(N__39981),
            .in2(_gnd_net_),
            .in3(N__39965),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_15_26_1  (
            .in0(N__40412),
            .in1(N__39951),
            .in2(_gnd_net_),
            .in3(N__39935),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_15_26_2  (
            .in0(N__40383),
            .in1(N__39919),
            .in2(_gnd_net_),
            .in3(N__39905),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_15_26_3  (
            .in0(N__40409),
            .in1(N__39894),
            .in2(_gnd_net_),
            .in3(N__39878),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_15_26_4  (
            .in0(N__40384),
            .in1(N__39873),
            .in2(_gnd_net_),
            .in3(N__39857),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_26_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_15_26_5  (
            .in0(N__40410),
            .in1(N__39852),
            .in2(_gnd_net_),
            .in3(N__39836),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_26_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_15_26_6  (
            .in0(N__40385),
            .in1(N__40251),
            .in2(_gnd_net_),
            .in3(N__40235),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_26_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_26_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_15_26_7  (
            .in0(N__40411),
            .in1(N__40219),
            .in2(_gnd_net_),
            .in3(N__40205),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__48334),
            .ce(N__40276),
            .sr(N__47861));
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_27_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_27_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_15_27_0  (
            .in0(N__40401),
            .in1(N__40194),
            .in2(_gnd_net_),
            .in3(N__40178),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_27_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_27_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_15_27_1  (
            .in0(N__40405),
            .in1(N__40167),
            .in2(_gnd_net_),
            .in3(N__40148),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_27_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_27_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_15_27_2  (
            .in0(N__40402),
            .in1(N__40132),
            .in2(_gnd_net_),
            .in3(N__40118),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_27_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_27_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_15_27_3  (
            .in0(N__40406),
            .in1(N__40102),
            .in2(_gnd_net_),
            .in3(N__40088),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_27_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_27_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_15_27_4  (
            .in0(N__40403),
            .in1(N__40083),
            .in2(_gnd_net_),
            .in3(N__40067),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_27_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_27_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_27_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_15_27_5  (
            .in0(N__40407),
            .in1(N__40057),
            .in2(_gnd_net_),
            .in3(N__40043),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_27_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_27_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_27_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_15_27_6  (
            .in0(N__40404),
            .in1(N__40597),
            .in2(_gnd_net_),
            .in3(N__40583),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_27_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_27_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_27_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_15_27_7  (
            .in0(N__40408),
            .in1(N__40572),
            .in2(_gnd_net_),
            .in3(N__40556),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__48333),
            .ce(N__40275),
            .sr(N__47868));
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_28_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_28_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_28_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_15_28_0  (
            .in0(N__40413),
            .in1(N__40545),
            .in2(_gnd_net_),
            .in3(N__40529),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_28_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__48331),
            .ce(N__40274),
            .sr(N__47872));
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_28_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_28_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_28_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_15_28_1  (
            .in0(N__40417),
            .in1(N__40518),
            .in2(_gnd_net_),
            .in3(N__40502),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__48331),
            .ce(N__40274),
            .sr(N__47872));
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_28_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_28_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_28_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_15_28_2  (
            .in0(N__40414),
            .in1(N__40486),
            .in2(_gnd_net_),
            .in3(N__40472),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__48331),
            .ce(N__40274),
            .sr(N__47872));
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_28_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_28_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_28_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_15_28_3  (
            .in0(N__40418),
            .in1(N__40456),
            .in2(_gnd_net_),
            .in3(N__40442),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__48331),
            .ce(N__40274),
            .sr(N__47872));
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_28_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_28_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_28_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_15_28_4  (
            .in0(N__40415),
            .in1(N__40435),
            .in2(_gnd_net_),
            .in3(N__40421),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__48331),
            .ce(N__40274),
            .sr(N__47872));
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_28_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_28_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_28_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_15_28_5  (
            .in0(N__40291),
            .in1(N__40416),
            .in2(_gnd_net_),
            .in3(N__40298),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48331),
            .ce(N__40274),
            .sr(N__47872));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_6_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_6_3  (
            .in0(N__41256),
            .in1(N__40764),
            .in2(N__41232),
            .in3(N__45595),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_6_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_6_4  (
            .in0(N__41280),
            .in1(N__40872),
            .in2(N__40850),
            .in3(N__40786),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_6_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_6_5  (
            .in0(N__41257),
            .in1(N__41281),
            .in2(N__41233),
            .in3(N__40873),
            .lcout(\delay_measurement_inst.N_265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_6_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_6_6  (
            .in0(_gnd_net_),
            .in1(N__40741),
            .in2(_gnd_net_),
            .in3(N__40717),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_287_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(N__45667),
            .in2(N__42544),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(N__45616),
            .in2(N__42520),
            .in3(N__40730),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__42942),
            .in2(N__42545),
            .in3(N__40706),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__42924),
            .in2(N__42521),
            .in3(N__40640),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__42943),
            .in2(N__42907),
            .in3(N__40613),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(N__42925),
            .in2(N__42883),
            .in3(N__41132),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(N__42860),
            .in2(N__42908),
            .in3(N__41081),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(N__42836),
            .in2(N__42884),
            .in3(N__41057),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48450),
            .ce(N__45564),
            .sr(N__47750));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__42859),
            .in2(N__42811),
            .in3(N__41036),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__42835),
            .in2(N__42787),
            .in3(N__41012),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__43125),
            .in2(N__42812),
            .in3(N__40988),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__43107),
            .in2(N__42788),
            .in3(N__40940),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__43126),
            .in2(N__43090),
            .in3(N__40883),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__43108),
            .in2(N__43066),
            .in3(N__40853),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__43043),
            .in2(N__43091),
            .in3(N__41264),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__43019),
            .in2(N__43067),
            .in3(N__41237),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48441),
            .ce(N__45565),
            .sr(N__47755));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__43042),
            .in2(N__42994),
            .in3(N__41204),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__43018),
            .in2(N__42970),
            .in3(N__41195),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__43320),
            .in2(N__42995),
            .in3(N__41186),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__43302),
            .in2(N__42971),
            .in3(N__41177),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__43321),
            .in2(N__43285),
            .in3(N__41165),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__43303),
            .in2(N__43261),
            .in3(N__41156),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__43238),
            .in2(N__43286),
            .in3(N__41513),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__43214),
            .in2(N__43262),
            .in3(N__41504),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48431),
            .ce(N__45567),
            .sr(N__47759));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__43237),
            .in2(N__43189),
            .in3(N__41489),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48423),
            .ce(N__45569),
            .sr(N__47769));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__43213),
            .in2(N__43165),
            .in3(N__41474),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48423),
            .ce(N__45569),
            .sr(N__47769));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__43141),
            .in2(N__43190),
            .in3(N__41459),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48423),
            .ce(N__45569),
            .sr(N__47769));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__43984),
            .in2(N__43166),
            .in3(N__41441),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48423),
            .ce(N__45569),
            .sr(N__47769));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41438),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48423),
            .ce(N__45569),
            .sr(N__47769));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_16_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_16_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__41342),
            .in2(N__41330),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_16_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_16_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__41306),
            .in2(_gnd_net_),
            .in3(N__41762),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_16_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__41759),
            .in2(N__41747),
            .in3(N__41717),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_16_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_16_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__41714),
            .in2(_gnd_net_),
            .in3(N__41687),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_16_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_16_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__41684),
            .in2(_gnd_net_),
            .in3(N__41657),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_16_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_16_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__41654),
            .in2(_gnd_net_),
            .in3(N__41624),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_16_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_16_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__41621),
            .in2(_gnd_net_),
            .in3(N__41588),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_16_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_16_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__41585),
            .in2(_gnd_net_),
            .in3(N__41549),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_16_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_16_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__41546),
            .in2(_gnd_net_),
            .in3(N__41522),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_16_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_16_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__41993),
            .in2(_gnd_net_),
            .in3(N__41963),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_16_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_16_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__41960),
            .in2(_gnd_net_),
            .in3(N__41930),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_16_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_16_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__41927),
            .in2(_gnd_net_),
            .in3(N__41897),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_16_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_16_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__41894),
            .in2(_gnd_net_),
            .in3(N__41864),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_16_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_16_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__41861),
            .in2(_gnd_net_),
            .in3(N__41831),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_16_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_16_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__41828),
            .in2(_gnd_net_),
            .in3(N__41798),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_16_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_16_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__43930),
            .in2(_gnd_net_),
            .in3(N__41795),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_16_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_16_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__41792),
            .in2(_gnd_net_),
            .in3(N__41774),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_16_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_16_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__42110),
            .in2(_gnd_net_),
            .in3(N__42092),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_16_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_16_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__42089),
            .in2(_gnd_net_),
            .in3(N__42077),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__42068),
            .in2(N__42044),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__46319),
            .in2(N__46354),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__42014),
            .in2(N__49349),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_16_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_16_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__49170),
            .in2(N__44138),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_16_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_16_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__44177),
            .in2(N__49350),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_16_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_16_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__49174),
            .in2(N__44219),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_16_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_16_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__41999),
            .in2(N__49351),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_16_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_16_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__49178),
            .in2(N__44276),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_16_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__49179),
            .in2(N__44591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_16_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__44423),
            .in2(N__49352),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_16_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__49183),
            .in2(N__42131),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_16_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__44486),
            .in2(N__49353),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_16_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__49187),
            .in2(N__44288),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_16_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__42122),
            .in2(N__49354),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_16_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__49191),
            .in2(N__44129),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_16_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__42116),
            .in2(N__49355),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_16_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__49068),
            .in2(N__44306),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_16_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__42380),
            .in2(N__49272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_16_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__49072),
            .in2(N__42317),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_16_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__44582),
            .in2(N__49273),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__49076),
            .in2(N__45359),
            .in3(N__42161),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(N__48782),
            .in2(N__49274),
            .in3(N__42152),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__49080),
            .in2(N__42341),
            .in3(N__42143),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(N__44294),
            .in2(N__49275),
            .in3(N__42134),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__42323),
            .in2(N__49276),
            .in3(N__42272),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__49087),
            .in2(N__42296),
            .in3(N__42263),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__42416),
            .in2(N__49277),
            .in3(N__42254),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__49091),
            .in2(N__42251),
            .in3(N__42227),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__47021),
            .in2(N__49278),
            .in3(N__42215),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__49095),
            .in2(N__45341),
            .in3(N__42203),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_16_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__42440),
            .in2(N__49279),
            .in3(N__42191),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_2_11_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_2_11_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_2_11_LC_16_17_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.control_input_RNO_2_11_LC_16_17_7  (
            .in0(N__49790),
            .in1(N__49099),
            .in2(_gnd_net_),
            .in3(N__42188),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_18_0  (
            .in0(N__49618),
            .in1(N__44205),
            .in2(N__49285),
            .in3(N__44757),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_18_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_18_1  (
            .in0(N__49106),
            .in1(N__49620),
            .in2(N__44378),
            .in3(N__44703),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_18_2  (
            .in0(N__49617),
            .in1(N__44262),
            .in2(N__49284),
            .in3(N__44817),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_3  (
            .in0(N__49103),
            .in1(N__49623),
            .in2(N__46931),
            .in3(N__46882),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_16_18_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_16_18_4  (
            .in0(N__49621),
            .in1(N__47437),
            .in2(N__49282),
            .in3(N__47386),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_5  (
            .in0(N__49104),
            .in1(N__49624),
            .in2(N__46550),
            .in3(N__46501),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_18_6  (
            .in0(N__49622),
            .in1(N__46855),
            .in2(N__49283),
            .in3(N__46810),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_18_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_18_7  (
            .in0(N__49105),
            .in1(N__49619),
            .in2(N__45191),
            .in3(N__44737),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_19_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_19_0  (
            .in0(N__49249),
            .in1(N__49757),
            .in2(N__46267),
            .in3(N__46219),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_16_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_16_19_1 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_16_19_1  (
            .in0(N__49754),
            .in1(N__46701),
            .in2(N__46648),
            .in3(N__49256),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_19_2 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_19_2  (
            .in0(N__49250),
            .in1(N__47356),
            .in2(N__47318),
            .in3(N__49756),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_19_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_19_3  (
            .in0(N__49753),
            .in1(N__49254),
            .in2(N__44576),
            .in3(N__44898),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_19_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_19_4  (
            .in0(N__44334),
            .in1(N__49751),
            .in2(N__49378),
            .in3(N__44976),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47426),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_19_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_19_6  (
            .in0(N__49248),
            .in1(N__49755),
            .in2(N__45287),
            .in3(N__45114),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_16_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_16_19_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_16_19_7  (
            .in0(N__49752),
            .in1(N__49255),
            .in2(N__46784),
            .in3(N__46732),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_20_0  (
            .in0(N__49763),
            .in1(N__47008),
            .in2(N__49379),
            .in3(N__46979),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_20_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_20_1  (
            .in0(N__49266),
            .in1(N__49762),
            .in2(N__46268),
            .in3(N__46218),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_20_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_20_2  (
            .in0(N__44193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_20_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_20_3  (
            .in0(N__47282),
            .in1(N__49761),
            .in2(N__49381),
            .in3(N__47255),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_4  (
            .in0(N__49765),
            .in1(N__47227),
            .in2(N__49380),
            .in3(N__47186),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44237),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_20_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_20_6  (
            .in0(N__49764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47159),
            .lcout(\current_shift_inst.un4_control_input_0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44151),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44355),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_16_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44317),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_2  (
            .in0(N__49785),
            .in1(N__47317),
            .in2(N__49433),
            .in3(N__47349),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44396),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_21_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_21_4  (
            .in0(N__46593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42477),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_6  (
            .in0(N__49786),
            .in1(N__47136),
            .in2(N__49432),
            .in3(N__47095),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46754),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48754),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_22_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__44507),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46904),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46832),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46238),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46990),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47336),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44556),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46521),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_24_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(N__47115),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_17_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_17_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_17_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42760),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48472),
            .ce(N__42710),
            .sr(N__47736));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_6_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_6_6  (
            .in0(N__42641),
            .in1(N__42620),
            .in2(_gnd_net_),
            .in3(N__42590),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_305_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0  (
            .in0(N__44113),
            .in1(N__45666),
            .in2(_gnd_net_),
            .in3(N__42551),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1  (
            .in0(N__44117),
            .in1(N__45615),
            .in2(_gnd_net_),
            .in3(N__42548),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2  (
            .in0(N__44114),
            .in1(N__42543),
            .in2(_gnd_net_),
            .in3(N__42524),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3  (
            .in0(N__44118),
            .in1(N__42519),
            .in2(_gnd_net_),
            .in3(N__42947),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4  (
            .in0(N__44115),
            .in1(N__42944),
            .in2(_gnd_net_),
            .in3(N__42929),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5  (
            .in0(N__44119),
            .in1(N__42926),
            .in2(_gnd_net_),
            .in3(N__42911),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6  (
            .in0(N__44116),
            .in1(N__42906),
            .in2(_gnd_net_),
            .in3(N__42887),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7  (
            .in0(N__44120),
            .in1(N__42882),
            .in2(_gnd_net_),
            .in3(N__42863),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__48461),
            .ce(N__43955),
            .sr(N__47742));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0  (
            .in0(N__44057),
            .in1(N__42858),
            .in2(_gnd_net_),
            .in3(N__42839),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1  (
            .in0(N__44080),
            .in1(N__42834),
            .in2(_gnd_net_),
            .in3(N__42815),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2  (
            .in0(N__44054),
            .in1(N__42810),
            .in2(_gnd_net_),
            .in3(N__42791),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3  (
            .in0(N__44077),
            .in1(N__42786),
            .in2(_gnd_net_),
            .in3(N__42767),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4  (
            .in0(N__44055),
            .in1(N__43127),
            .in2(_gnd_net_),
            .in3(N__43112),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5  (
            .in0(N__44078),
            .in1(N__43109),
            .in2(_gnd_net_),
            .in3(N__43094),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6  (
            .in0(N__44056),
            .in1(N__43089),
            .in2(_gnd_net_),
            .in3(N__43070),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7  (
            .in0(N__44079),
            .in1(N__43065),
            .in2(_gnd_net_),
            .in3(N__43046),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__48451),
            .ce(N__43965),
            .sr(N__47751));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0  (
            .in0(N__44091),
            .in1(N__43041),
            .in2(_gnd_net_),
            .in3(N__43022),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1  (
            .in0(N__44085),
            .in1(N__43017),
            .in2(_gnd_net_),
            .in3(N__42998),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2  (
            .in0(N__44092),
            .in1(N__42993),
            .in2(_gnd_net_),
            .in3(N__42974),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3  (
            .in0(N__44086),
            .in1(N__42969),
            .in2(_gnd_net_),
            .in3(N__42950),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4  (
            .in0(N__44093),
            .in1(N__43322),
            .in2(_gnd_net_),
            .in3(N__43307),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5  (
            .in0(N__44087),
            .in1(N__43304),
            .in2(_gnd_net_),
            .in3(N__43289),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6  (
            .in0(N__44094),
            .in1(N__43284),
            .in2(_gnd_net_),
            .in3(N__43265),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7  (
            .in0(N__44088),
            .in1(N__43260),
            .in2(_gnd_net_),
            .in3(N__43241),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__48442),
            .ce(N__43973),
            .sr(N__47756));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0  (
            .in0(N__44081),
            .in1(N__43236),
            .in2(_gnd_net_),
            .in3(N__43217),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__48432),
            .ce(N__43969),
            .sr(N__47760));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1  (
            .in0(N__44089),
            .in1(N__43212),
            .in2(_gnd_net_),
            .in3(N__43193),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__48432),
            .ce(N__43969),
            .sr(N__47760));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2  (
            .in0(N__44082),
            .in1(N__43188),
            .in2(_gnd_net_),
            .in3(N__43169),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__48432),
            .ce(N__43969),
            .sr(N__47760));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3  (
            .in0(N__44090),
            .in1(N__43164),
            .in2(_gnd_net_),
            .in3(N__43145),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__48432),
            .ce(N__43969),
            .sr(N__47760));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4  (
            .in0(N__44083),
            .in1(N__43142),
            .in2(_gnd_net_),
            .in3(N__43130),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__48432),
            .ce(N__43969),
            .sr(N__47760));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5  (
            .in0(N__43985),
            .in1(N__44084),
            .in2(_gnd_net_),
            .in3(N__43988),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48432),
            .ce(N__43969),
            .sr(N__47760));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_0  (
            .in0(N__43561),
            .in1(N__43826),
            .in2(N__43683),
            .in3(N__43937),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48424),
            .ce(),
            .sr(N__47770));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_11_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__43559),
            .in2(_gnd_net_),
            .in3(N__43824),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_11_3 .LUT_INIT=16'b1010100010111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_17_11_3  (
            .in0(N__43402),
            .in1(N__43448),
            .in2(N__43892),
            .in3(N__43889),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48424),
            .ce(),
            .sr(N__47770));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__43401),
            .in2(_gnd_net_),
            .in3(N__43333),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_11_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_11_7  (
            .in0(N__43825),
            .in1(N__43640),
            .in2(_gnd_net_),
            .in3(N__43560),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_17_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_17_12_6 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_0_LC_17_12_6  (
            .in0(N__43435),
            .in1(N__43403),
            .in2(N__43388),
            .in3(N__43334),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48412),
            .ce(),
            .sr(N__47773));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_13_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_13_2  (
            .in0(N__48687),
            .in1(N__44263),
            .in2(_gnd_net_),
            .in3(N__44821),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_14_0 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_14_0  (
            .in0(N__44759),
            .in1(N__49748),
            .in2(N__44210),
            .in3(N__49443),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_14_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_14_1  (
            .in0(N__49747),
            .in1(N__49427),
            .in2(N__44267),
            .in3(N__44822),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2  (
            .in0(N__48670),
            .in1(N__46612),
            .in2(_gnd_net_),
            .in3(N__46579),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3  (
            .in0(N__48689),
            .in1(N__44206),
            .in2(_gnd_net_),
            .in3(N__44758),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_17_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_17_14_4  (
            .in0(N__49746),
            .in1(N__46613),
            .in2(N__49450),
            .in3(N__46580),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5  (
            .in0(N__48688),
            .in1(N__45236),
            .in2(_gnd_net_),
            .in3(N__44788),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6  (
            .in0(N__48669),
            .in1(N__44167),
            .in2(_gnd_net_),
            .in3(N__44460),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_14_7 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_14_7  (
            .in0(N__44461),
            .in1(N__49745),
            .in2(N__44171),
            .in3(N__49423),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_15_0 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_15_0  (
            .in0(N__44978),
            .in1(N__49776),
            .in2(N__44339),
            .in3(N__49439),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_15_1  (
            .in0(N__49775),
            .in1(N__44377),
            .in2(N__49454),
            .in3(N__44705),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_2  (
            .in0(N__44417),
            .in1(N__48673),
            .in2(_gnd_net_),
            .in3(N__44664),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3  (
            .in0(N__48672),
            .in1(N__44376),
            .in2(_gnd_net_),
            .in3(N__44704),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_4  (
            .in0(N__47068),
            .in1(N__48676),
            .in2(_gnd_net_),
            .in3(N__44943),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_5  (
            .in0(N__48675),
            .in1(N__44335),
            .in2(_gnd_net_),
            .in3(N__44977),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6  (
            .in0(N__44535),
            .in1(N__48674),
            .in2(_gnd_net_),
            .in3(N__44622),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_15_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_15_7  (
            .in0(N__48671),
            .in1(N__45189),
            .in2(_gnd_net_),
            .in3(N__44738),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_17_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_17_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_17_16_0  (
            .in0(N__44572),
            .in1(N__49780),
            .in2(N__49457),
            .in3(N__44902),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_16_1  (
            .in0(N__49782),
            .in1(N__45283),
            .in2(N__49434),
            .in3(N__45116),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_16_2 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_16_2  (
            .in0(N__47390),
            .in1(N__49779),
            .in2(N__47438),
            .in3(N__49401),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_16_3  (
            .in0(N__49777),
            .in1(N__45190),
            .in2(N__49435),
            .in3(N__44736),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_17_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_17_16_4 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_17_16_4  (
            .in0(N__46649),
            .in1(N__49781),
            .in2(N__46706),
            .in3(N__49402),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_5  (
            .in0(N__48665),
            .in1(_gnd_net_),
            .in2(N__44903),
            .in3(N__44571),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_16_6 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_16_6  (
            .in0(N__44626),
            .in1(N__49778),
            .in2(N__44540),
            .in3(N__49400),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_7  (
            .in0(N__48666),
            .in1(N__45282),
            .in2(_gnd_net_),
            .in3(N__45115),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__46361),
            .in2(N__45326),
            .in3(N__45324),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__46937),
            .in2(_gnd_net_),
            .in3(N__44480),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__44477),
            .in2(_gnd_net_),
            .in3(N__44441),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__44438),
            .in2(_gnd_net_),
            .in3(N__44426),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__44831),
            .in2(_gnd_net_),
            .in3(N__44798),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__45200),
            .in2(_gnd_net_),
            .in3(N__44771),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__44768),
            .in2(_gnd_net_),
            .in3(N__44741),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__45149),
            .in2(_gnd_net_),
            .in3(N__44717),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__44714),
            .in2(_gnd_net_),
            .in3(N__44687),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__44684),
            .in2(_gnd_net_),
            .in3(N__44642),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__44639),
            .in2(_gnd_net_),
            .in3(N__44603),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__44600),
            .in2(_gnd_net_),
            .in3(N__44594),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__45029),
            .in2(_gnd_net_),
            .in3(N__44993),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__44990),
            .in2(_gnd_net_),
            .in3(N__44960),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__47027),
            .in2(_gnd_net_),
            .in3(N__44918),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__44915),
            .in2(_gnd_net_),
            .in3(N__44882),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__44879),
            .in2(_gnd_net_),
            .in3(N__44870),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__44867),
            .in2(_gnd_net_),
            .in3(N__44855),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__44852),
            .in2(_gnd_net_),
            .in3(N__44837),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__46475),
            .in2(_gnd_net_),
            .in3(N__44834),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__45140),
            .in2(_gnd_net_),
            .in3(N__45131),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__45128),
            .in2(_gnd_net_),
            .in3(N__45119),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__45245),
            .in2(_gnd_net_),
            .in3(N__45098),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__45095),
            .in2(_gnd_net_),
            .in3(N__45083),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__45080),
            .in2(_gnd_net_),
            .in3(N__45071),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__45068),
            .in2(_gnd_net_),
            .in3(N__45059),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__45056),
            .in2(_gnd_net_),
            .in3(N__45044),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__45041),
            .in2(_gnd_net_),
            .in3(N__45032),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__45677),
            .in2(_gnd_net_),
            .in3(N__45365),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45362),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_20_6  (
            .in0(N__49784),
            .in1(N__47288),
            .in2(N__49431),
            .in3(N__47254),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_17_20_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_17_20_7  (
            .in0(N__49766),
            .in1(N__49377),
            .in2(N__47228),
            .in3(N__47185),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48495),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_21_3 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_21_3  (
            .in0(N__48496),
            .in1(_gnd_net_),
            .in2(N__45290),
            .in3(N__48575),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45281),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45227),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45171),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47205),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45668),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48473),
            .ce(N__45566),
            .sr(N__47737));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45617),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48468),
            .ce(N__45568),
            .sr(N__47739));
    defparam \phase_controller_inst1.state_4_LC_18_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_18_11_2 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_18_11_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__45510),
            .in2(_gnd_net_),
            .in3(N__45458),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48433),
            .ce(),
            .sr(N__47761));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_18_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_18_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__45433),
            .in2(N__45404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_18_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_18_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__46277),
            .in2(N__46148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_18_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_18_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__46172),
            .in2(N__46116),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_18_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_18_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__45377),
            .in2(N__46149),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_18_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_18_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__45371),
            .in2(N__46117),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_18_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_18_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__45722),
            .in2(N__46150),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_18_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_18_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__45716),
            .in2(N__46118),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_18_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_18_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__45710),
            .in2(N__46151),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_18_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_18_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__46129),
            .in2(N__45704),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_18_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_18_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__45695),
            .in2(N__46147),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_18_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_18_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__45689),
            .in2(N__46113),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_18_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_18_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__45683),
            .in2(N__46145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_18_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_18_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__47369),
            .in2(N__46114),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_18_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_18_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__46068),
            .in2(N__45752),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_18_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_18_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__45740),
            .in2(N__46115),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_18_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_18_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__45734),
            .in2(N__46146),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_18_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_18_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__45728),
            .in2(N__46119),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_18_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_18_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__46715),
            .in2(N__46059),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_18_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_18_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__46793),
            .in2(N__46120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_18_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_18_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__46622),
            .in2(N__46060),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_18_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_18_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__47237),
            .in2(N__46121),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_18_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_18_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__48731),
            .in2(N__46061),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_18_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_18_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__46865),
            .in2(N__46122),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_18_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_18_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__46094),
            .in2(N__46160),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_18_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_18_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__46484),
            .in2(N__46035),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_18_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_18_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__46199),
            .in2(N__46039),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_18_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_18_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__47297),
            .in2(N__46036),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_18_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_18_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__47078),
            .in2(N__46040),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_18_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_18_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__49820),
            .in2(N__46037),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_18_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_18_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__47168),
            .in2(N__46041),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_18_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_18_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__47147),
            .in2(N__46038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_16_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__49783),
            .in2(_gnd_net_),
            .in3(N__46469),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_17_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_17_0  (
            .in0(N__49707),
            .in1(N__46303),
            .in2(N__46355),
            .in3(N__46291),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46394),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48390),
            .ce(N__48017),
            .sr(N__47790));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46289),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_17_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_17_3  (
            .in0(N__46292),
            .in1(N__49708),
            .in2(N__46307),
            .in3(N__46353),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_17_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_17_4  (
            .in0(N__48604),
            .in1(N__46302),
            .in2(_gnd_net_),
            .in3(N__46290),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_17_7  (
            .in0(N__49709),
            .in1(N__46266),
            .in2(_gnd_net_),
            .in3(N__46220),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_18_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_18_0  (
            .in0(N__46964),
            .in1(N__48605),
            .in2(_gnd_net_),
            .in3(N__46183),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46963),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_18_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_18_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_18_18_2  (
            .in0(N__48668),
            .in1(N__46930),
            .in2(_gnd_net_),
            .in3(N__46881),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_18_3  (
            .in0(N__48606),
            .in1(N__46856),
            .in2(_gnd_net_),
            .in3(N__46809),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_18_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_18_4  (
            .in0(N__48667),
            .in1(N__46782),
            .in2(_gnd_net_),
            .in3(N__46731),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_18_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_18_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_18_18_5  (
            .in0(N__48607),
            .in1(N__46702),
            .in2(_gnd_net_),
            .in3(N__46638),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_18_6  (
            .in0(N__49710),
            .in1(N__46611),
            .in2(N__49455),
            .in3(N__46578),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_18_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_18_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_18_18_7  (
            .in0(N__48608),
            .in1(N__46546),
            .in2(_gnd_net_),
            .in3(N__46500),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47286),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_19_1  (
            .in0(N__48658),
            .in1(N__47427),
            .in2(_gnd_net_),
            .in3(N__47385),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_18_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_18_19_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_18_19_2  (
            .in0(N__49738),
            .in1(N__47357),
            .in2(_gnd_net_),
            .in3(N__47313),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_19_3 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_19_3  (
            .in0(N__47287),
            .in1(_gnd_net_),
            .in2(N__48685),
            .in3(N__47253),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_18_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_18_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_18_19_4  (
            .in0(N__49739),
            .in1(N__47223),
            .in2(_gnd_net_),
            .in3(N__47184),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_19_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__49740),
            .in2(_gnd_net_),
            .in3(N__47158),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_18_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_18_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_18_19_6  (
            .in0(N__49737),
            .in1(N__47138),
            .in2(_gnd_net_),
            .in3(N__47094),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47067),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_18_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_18_20_1 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_18_20_1  (
            .in0(N__46978),
            .in1(N__49735),
            .in2(N__47009),
            .in3(N__49370),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_18_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_18_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_18_20_2  (
            .in0(N__49733),
            .in1(N__47004),
            .in2(_gnd_net_),
            .in3(N__46977),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_1_11_LC_18_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_1_11_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_1_11_LC_18_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_RNO_1_11_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__49736),
            .in2(_gnd_net_),
            .in3(N__49369),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_20_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_20_4  (
            .in0(N__49732),
            .in1(N__48769),
            .in2(N__49430),
            .in3(N__48742),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_20_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_20_5  (
            .in0(N__48743),
            .in1(N__49734),
            .in2(N__49456),
            .in3(N__48770),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_18_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_18_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_18_20_6  (
            .in0(N__48603),
            .in1(N__48768),
            .in2(_gnd_net_),
            .in3(N__48741),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48721),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48375),
            .ce(N__48012),
            .sr(N__47802));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48544),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48370),
            .ce(N__48016),
            .sr(N__47806));
endmodule // MAIN
