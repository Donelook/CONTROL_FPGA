// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 24 2025 22:26:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__48680;
    wire N__48679;
    wire N__48678;
    wire N__48669;
    wire N__48668;
    wire N__48667;
    wire N__48660;
    wire N__48659;
    wire N__48658;
    wire N__48651;
    wire N__48650;
    wire N__48649;
    wire N__48642;
    wire N__48641;
    wire N__48640;
    wire N__48633;
    wire N__48632;
    wire N__48631;
    wire N__48624;
    wire N__48623;
    wire N__48622;
    wire N__48615;
    wire N__48614;
    wire N__48613;
    wire N__48606;
    wire N__48605;
    wire N__48604;
    wire N__48597;
    wire N__48596;
    wire N__48595;
    wire N__48588;
    wire N__48587;
    wire N__48586;
    wire N__48579;
    wire N__48578;
    wire N__48577;
    wire N__48570;
    wire N__48569;
    wire N__48568;
    wire N__48551;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48543;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48529;
    wire N__48524;
    wire N__48521;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48509;
    wire N__48506;
    wire N__48505;
    wire N__48504;
    wire N__48499;
    wire N__48496;
    wire N__48495;
    wire N__48494;
    wire N__48491;
    wire N__48488;
    wire N__48485;
    wire N__48482;
    wire N__48479;
    wire N__48472;
    wire N__48467;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48459;
    wire N__48454;
    wire N__48451;
    wire N__48446;
    wire N__48443;
    wire N__48442;
    wire N__48439;
    wire N__48438;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48417;
    wire N__48410;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48402;
    wire N__48397;
    wire N__48394;
    wire N__48389;
    wire N__48388;
    wire N__48385;
    wire N__48382;
    wire N__48377;
    wire N__48374;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48366;
    wire N__48361;
    wire N__48358;
    wire N__48357;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48338;
    wire N__48335;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48327;
    wire N__48322;
    wire N__48319;
    wire N__48318;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48290;
    wire N__48287;
    wire N__48284;
    wire N__48283;
    wire N__48282;
    wire N__48281;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48275;
    wire N__48274;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48262;
    wire N__48261;
    wire N__48260;
    wire N__48259;
    wire N__48258;
    wire N__48257;
    wire N__48254;
    wire N__48253;
    wire N__48252;
    wire N__48247;
    wire N__48240;
    wire N__48231;
    wire N__48228;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48216;
    wire N__48215;
    wire N__48212;
    wire N__48211;
    wire N__48208;
    wire N__48203;
    wire N__48196;
    wire N__48191;
    wire N__48178;
    wire N__48173;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48155;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48133;
    wire N__48130;
    wire N__48125;
    wire N__48122;
    wire N__48121;
    wire N__48120;
    wire N__48119;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48107;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48092;
    wire N__48091;
    wire N__48090;
    wire N__48081;
    wire N__48080;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48059;
    wire N__48056;
    wire N__48055;
    wire N__48054;
    wire N__48051;
    wire N__48048;
    wire N__48045;
    wire N__48044;
    wire N__48041;
    wire N__48038;
    wire N__48035;
    wire N__48032;
    wire N__48027;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48013;
    wire N__48008;
    wire N__48007;
    wire N__48006;
    wire N__48005;
    wire N__48004;
    wire N__48003;
    wire N__48002;
    wire N__48001;
    wire N__48000;
    wire N__47999;
    wire N__47998;
    wire N__47997;
    wire N__47996;
    wire N__47995;
    wire N__47994;
    wire N__47993;
    wire N__47992;
    wire N__47991;
    wire N__47990;
    wire N__47989;
    wire N__47988;
    wire N__47987;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47983;
    wire N__47982;
    wire N__47981;
    wire N__47980;
    wire N__47979;
    wire N__47978;
    wire N__47977;
    wire N__47976;
    wire N__47975;
    wire N__47974;
    wire N__47973;
    wire N__47972;
    wire N__47971;
    wire N__47970;
    wire N__47969;
    wire N__47968;
    wire N__47967;
    wire N__47966;
    wire N__47965;
    wire N__47964;
    wire N__47963;
    wire N__47962;
    wire N__47961;
    wire N__47960;
    wire N__47959;
    wire N__47958;
    wire N__47957;
    wire N__47956;
    wire N__47955;
    wire N__47954;
    wire N__47953;
    wire N__47952;
    wire N__47951;
    wire N__47950;
    wire N__47949;
    wire N__47948;
    wire N__47947;
    wire N__47946;
    wire N__47945;
    wire N__47944;
    wire N__47943;
    wire N__47942;
    wire N__47941;
    wire N__47940;
    wire N__47939;
    wire N__47938;
    wire N__47937;
    wire N__47936;
    wire N__47935;
    wire N__47934;
    wire N__47933;
    wire N__47932;
    wire N__47931;
    wire N__47930;
    wire N__47929;
    wire N__47928;
    wire N__47927;
    wire N__47926;
    wire N__47925;
    wire N__47924;
    wire N__47923;
    wire N__47922;
    wire N__47921;
    wire N__47920;
    wire N__47919;
    wire N__47918;
    wire N__47917;
    wire N__47916;
    wire N__47915;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47911;
    wire N__47910;
    wire N__47909;
    wire N__47908;
    wire N__47907;
    wire N__47906;
    wire N__47905;
    wire N__47904;
    wire N__47903;
    wire N__47902;
    wire N__47901;
    wire N__47900;
    wire N__47899;
    wire N__47898;
    wire N__47897;
    wire N__47896;
    wire N__47895;
    wire N__47894;
    wire N__47893;
    wire N__47892;
    wire N__47891;
    wire N__47890;
    wire N__47889;
    wire N__47888;
    wire N__47887;
    wire N__47886;
    wire N__47885;
    wire N__47884;
    wire N__47883;
    wire N__47882;
    wire N__47881;
    wire N__47880;
    wire N__47879;
    wire N__47878;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47860;
    wire N__47859;
    wire N__47858;
    wire N__47857;
    wire N__47856;
    wire N__47855;
    wire N__47854;
    wire N__47853;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47522;
    wire N__47519;
    wire N__47518;
    wire N__47515;
    wire N__47512;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47492;
    wire N__47491;
    wire N__47490;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47465;
    wire N__47464;
    wire N__47463;
    wire N__47462;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47438;
    wire N__47435;
    wire N__47432;
    wire N__47429;
    wire N__47426;
    wire N__47423;
    wire N__47422;
    wire N__47421;
    wire N__47418;
    wire N__47417;
    wire N__47416;
    wire N__47415;
    wire N__47414;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47408;
    wire N__47407;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47403;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47398;
    wire N__47397;
    wire N__47396;
    wire N__47395;
    wire N__47394;
    wire N__47393;
    wire N__47392;
    wire N__47391;
    wire N__47390;
    wire N__47389;
    wire N__47388;
    wire N__47387;
    wire N__47386;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47374;
    wire N__47373;
    wire N__47372;
    wire N__47371;
    wire N__47370;
    wire N__47369;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47355;
    wire N__47354;
    wire N__47353;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47332;
    wire N__47331;
    wire N__47330;
    wire N__47329;
    wire N__47328;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47309;
    wire N__47308;
    wire N__47307;
    wire N__47306;
    wire N__47305;
    wire N__47304;
    wire N__47303;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47299;
    wire N__47298;
    wire N__47297;
    wire N__47296;
    wire N__47295;
    wire N__47294;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47290;
    wire N__47289;
    wire N__47288;
    wire N__47287;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47279;
    wire N__47278;
    wire N__47277;
    wire N__47276;
    wire N__47275;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__46979;
    wire N__46976;
    wire N__46973;
    wire N__46970;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46946;
    wire N__46945;
    wire N__46942;
    wire N__46941;
    wire N__46938;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46924;
    wire N__46919;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46911;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46897;
    wire N__46894;
    wire N__46889;
    wire N__46888;
    wire N__46885;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46850;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46823;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46815;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46803;
    wire N__46798;
    wire N__46795;
    wire N__46792;
    wire N__46787;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46777;
    wire N__46774;
    wire N__46771;
    wire N__46768;
    wire N__46763;
    wire N__46760;
    wire N__46759;
    wire N__46758;
    wire N__46755;
    wire N__46752;
    wire N__46749;
    wire N__46742;
    wire N__46739;
    wire N__46736;
    wire N__46735;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46719;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46700;
    wire N__46699;
    wire N__46696;
    wire N__46693;
    wire N__46690;
    wire N__46687;
    wire N__46682;
    wire N__46679;
    wire N__46678;
    wire N__46675;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46665;
    wire N__46662;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46648;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46637;
    wire N__46630;
    wire N__46627;
    wire N__46622;
    wire N__46619;
    wire N__46616;
    wire N__46615;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46598;
    wire N__46595;
    wire N__46592;
    wire N__46591;
    wire N__46588;
    wire N__46585;
    wire N__46582;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46568;
    wire N__46565;
    wire N__46564;
    wire N__46563;
    wire N__46560;
    wire N__46557;
    wire N__46554;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46540;
    wire N__46539;
    wire N__46538;
    wire N__46537;
    wire N__46536;
    wire N__46535;
    wire N__46534;
    wire N__46525;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46499;
    wire N__46498;
    wire N__46497;
    wire N__46490;
    wire N__46489;
    wire N__46488;
    wire N__46487;
    wire N__46484;
    wire N__46477;
    wire N__46472;
    wire N__46469;
    wire N__46468;
    wire N__46467;
    wire N__46464;
    wire N__46461;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46449;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46433;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46394;
    wire N__46391;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46364;
    wire N__46363;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46349;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46341;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46329;
    wire N__46322;
    wire N__46319;
    wire N__46318;
    wire N__46317;
    wire N__46314;
    wire N__46313;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46298;
    wire N__46295;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46277;
    wire N__46276;
    wire N__46275;
    wire N__46274;
    wire N__46273;
    wire N__46272;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46260;
    wire N__46255;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46226;
    wire N__46217;
    wire N__46214;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46206;
    wire N__46205;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46191;
    wire N__46184;
    wire N__46183;
    wire N__46182;
    wire N__46181;
    wire N__46180;
    wire N__46179;
    wire N__46178;
    wire N__46177;
    wire N__46174;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46156;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46132;
    wire N__46127;
    wire N__46120;
    wire N__46115;
    wire N__46110;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46091;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46067;
    wire N__46064;
    wire N__46061;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46048;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46028;
    wire N__46025;
    wire N__46022;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46009;
    wire N__46006;
    wire N__46003;
    wire N__46000;
    wire N__45993;
    wire N__45986;
    wire N__45983;
    wire N__45980;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45953;
    wire N__45950;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45940;
    wire N__45937;
    wire N__45934;
    wire N__45931;
    wire N__45926;
    wire N__45925;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45878;
    wire N__45875;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45832;
    wire N__45829;
    wire N__45826;
    wire N__45823;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45806;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45778;
    wire N__45775;
    wire N__45772;
    wire N__45769;
    wire N__45764;
    wire N__45761;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45728;
    wire N__45725;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45713;
    wire N__45712;
    wire N__45709;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45693;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45568;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45521;
    wire N__45518;
    wire N__45515;
    wire N__45514;
    wire N__45511;
    wire N__45508;
    wire N__45505;
    wire N__45500;
    wire N__45497;
    wire N__45494;
    wire N__45491;
    wire N__45488;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45446;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45436;
    wire N__45435;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45419;
    wire N__45416;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45406;
    wire N__45401;
    wire N__45398;
    wire N__45395;
    wire N__45392;
    wire N__45389;
    wire N__45388;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45377;
    wire N__45374;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45328;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45310;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45295;
    wire N__45292;
    wire N__45289;
    wire N__45284;
    wire N__45281;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45254;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45230;
    wire N__45227;
    wire N__45224;
    wire N__45221;
    wire N__45220;
    wire N__45217;
    wire N__45214;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45188;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45167;
    wire N__45164;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45140;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45132;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45106;
    wire N__45101;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45066;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45027;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__45001;
    wire N__45000;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44971;
    wire N__44968;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44948;
    wire N__44945;
    wire N__44942;
    wire N__44939;
    wire N__44936;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44909;
    wire N__44906;
    wire N__44903;
    wire N__44900;
    wire N__44897;
    wire N__44894;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44879;
    wire N__44878;
    wire N__44875;
    wire N__44872;
    wire N__44871;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44855;
    wire N__44852;
    wire N__44849;
    wire N__44846;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44835;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44819;
    wire N__44816;
    wire N__44815;
    wire N__44812;
    wire N__44809;
    wire N__44808;
    wire N__44803;
    wire N__44800;
    wire N__44797;
    wire N__44792;
    wire N__44789;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44781;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44765;
    wire N__44762;
    wire N__44761;
    wire N__44760;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44744;
    wire N__44741;
    wire N__44740;
    wire N__44739;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44723;
    wire N__44720;
    wire N__44719;
    wire N__44716;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44701;
    wire N__44696;
    wire N__44693;
    wire N__44692;
    wire N__44689;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44669;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44659;
    wire N__44656;
    wire N__44653;
    wire N__44652;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44636;
    wire N__44633;
    wire N__44630;
    wire N__44627;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44619;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44603;
    wire N__44600;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44592;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44576;
    wire N__44573;
    wire N__44572;
    wire N__44567;
    wire N__44566;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44552;
    wire N__44549;
    wire N__44548;
    wire N__44543;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44528;
    wire N__44525;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44514;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44498;
    wire N__44495;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44483;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44461;
    wire N__44458;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44431;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44414;
    wire N__44411;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44400;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44384;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44374;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44357;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44341;
    wire N__44336;
    wire N__44333;
    wire N__44332;
    wire N__44331;
    wire N__44330;
    wire N__44329;
    wire N__44328;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44298;
    wire N__44293;
    wire N__44290;
    wire N__44285;
    wire N__44284;
    wire N__44281;
    wire N__44278;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44261;
    wire N__44258;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44236;
    wire N__44233;
    wire N__44228;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44204;
    wire N__44201;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44189;
    wire N__44186;
    wire N__44185;
    wire N__44184;
    wire N__44183;
    wire N__44182;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44168;
    wire N__44165;
    wire N__44156;
    wire N__44153;
    wire N__44150;
    wire N__44149;
    wire N__44146;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44138;
    wire N__44135;
    wire N__44134;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44107;
    wire N__44102;
    wire N__44099;
    wire N__44090;
    wire N__44087;
    wire N__44084;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44071;
    wire N__44068;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44032;
    wire N__44021;
    wire N__44020;
    wire N__44017;
    wire N__44016;
    wire N__44015;
    wire N__44014;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43977;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43956;
    wire N__43951;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43943;
    wire N__43940;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43928;
    wire N__43925;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43900;
    wire N__43897;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43880;
    wire N__43879;
    wire N__43876;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43859;
    wire N__43856;
    wire N__43855;
    wire N__43854;
    wire N__43853;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43845;
    wire N__43844;
    wire N__43843;
    wire N__43842;
    wire N__43841;
    wire N__43840;
    wire N__43839;
    wire N__43836;
    wire N__43835;
    wire N__43834;
    wire N__43833;
    wire N__43830;
    wire N__43829;
    wire N__43828;
    wire N__43827;
    wire N__43826;
    wire N__43825;
    wire N__43824;
    wire N__43823;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43799;
    wire N__43796;
    wire N__43791;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43767;
    wire N__43764;
    wire N__43755;
    wire N__43750;
    wire N__43747;
    wire N__43740;
    wire N__43733;
    wire N__43732;
    wire N__43729;
    wire N__43728;
    wire N__43725;
    wire N__43724;
    wire N__43723;
    wire N__43722;
    wire N__43721;
    wire N__43720;
    wire N__43715;
    wire N__43714;
    wire N__43713;
    wire N__43712;
    wire N__43711;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43703;
    wire N__43702;
    wire N__43701;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43668;
    wire N__43667;
    wire N__43666;
    wire N__43665;
    wire N__43664;
    wire N__43661;
    wire N__43660;
    wire N__43657;
    wire N__43640;
    wire N__43635;
    wire N__43618;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43600;
    wire N__43589;
    wire N__43588;
    wire N__43587;
    wire N__43586;
    wire N__43585;
    wire N__43584;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43571;
    wire N__43570;
    wire N__43569;
    wire N__43568;
    wire N__43565;
    wire N__43564;
    wire N__43561;
    wire N__43560;
    wire N__43559;
    wire N__43558;
    wire N__43557;
    wire N__43556;
    wire N__43555;
    wire N__43554;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43540;
    wire N__43529;
    wire N__43526;
    wire N__43521;
    wire N__43520;
    wire N__43519;
    wire N__43516;
    wire N__43499;
    wire N__43494;
    wire N__43485;
    wire N__43480;
    wire N__43477;
    wire N__43470;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43445;
    wire N__43442;
    wire N__43441;
    wire N__43440;
    wire N__43439;
    wire N__43438;
    wire N__43437;
    wire N__43436;
    wire N__43435;
    wire N__43434;
    wire N__43431;
    wire N__43424;
    wire N__43413;
    wire N__43412;
    wire N__43411;
    wire N__43410;
    wire N__43409;
    wire N__43408;
    wire N__43407;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43382;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43354;
    wire N__43353;
    wire N__43352;
    wire N__43349;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43325;
    wire N__43318;
    wire N__43315;
    wire N__43310;
    wire N__43309;
    wire N__43304;
    wire N__43303;
    wire N__43302;
    wire N__43301;
    wire N__43300;
    wire N__43299;
    wire N__43298;
    wire N__43297;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43281;
    wire N__43274;
    wire N__43265;
    wire N__43264;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43249;
    wire N__43244;
    wire N__43243;
    wire N__43238;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43228;
    wire N__43223;
    wire N__43222;
    wire N__43219;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43190;
    wire N__43189;
    wire N__43188;
    wire N__43187;
    wire N__43186;
    wire N__43185;
    wire N__43176;
    wire N__43171;
    wire N__43166;
    wire N__43165;
    wire N__43164;
    wire N__43163;
    wire N__43162;
    wire N__43161;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43143;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43127;
    wire N__43124;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43112;
    wire N__43111;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43103;
    wire N__43100;
    wire N__43095;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43071;
    wire N__43064;
    wire N__43063;
    wire N__43062;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43050;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43033;
    wire N__43032;
    wire N__43029;
    wire N__43024;
    wire N__43023;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43015;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42989;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42981;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42905;
    wire N__42904;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42894;
    wire N__42893;
    wire N__42892;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42877;
    wire N__42874;
    wire N__42863;
    wire N__42862;
    wire N__42861;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42827;
    wire N__42824;
    wire N__42823;
    wire N__42818;
    wire N__42817;
    wire N__42814;
    wire N__42813;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42785;
    wire N__42782;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42774;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42739;
    wire N__42738;
    wire N__42737;
    wire N__42736;
    wire N__42735;
    wire N__42734;
    wire N__42733;
    wire N__42724;
    wire N__42723;
    wire N__42722;
    wire N__42721;
    wire N__42720;
    wire N__42719;
    wire N__42718;
    wire N__42717;
    wire N__42716;
    wire N__42715;
    wire N__42714;
    wire N__42713;
    wire N__42712;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42706;
    wire N__42705;
    wire N__42704;
    wire N__42703;
    wire N__42702;
    wire N__42693;
    wire N__42690;
    wire N__42681;
    wire N__42672;
    wire N__42663;
    wire N__42654;
    wire N__42649;
    wire N__42640;
    wire N__42633;
    wire N__42626;
    wire N__42621;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42602;
    wire N__42599;
    wire N__42596;
    wire N__42595;
    wire N__42592;
    wire N__42591;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42557;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42533;
    wire N__42530;
    wire N__42527;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42506;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42476;
    wire N__42475;
    wire N__42474;
    wire N__42471;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42437;
    wire N__42436;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42409;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42395;
    wire N__42392;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42380;
    wire N__42379;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42338;
    wire N__42335;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42319;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42289;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42269;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42259;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42229;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42199;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42170;
    wire N__42169;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42139;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42119;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42104;
    wire N__42101;
    wire N__42098;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42074;
    wire N__42073;
    wire N__42070;
    wire N__42067;
    wire N__42064;
    wire N__42059;
    wire N__42056;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42046;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42026;
    wire N__42023;
    wire N__42020;
    wire N__42017;
    wire N__42016;
    wire N__42013;
    wire N__42012;
    wire N__42011;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41987;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41970;
    wire N__41963;
    wire N__41960;
    wire N__41959;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41939;
    wire N__41936;
    wire N__41935;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41915;
    wire N__41912;
    wire N__41911;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41867;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41801;
    wire N__41798;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41780;
    wire N__41777;
    wire N__41776;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41756;
    wire N__41753;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41735;
    wire N__41732;
    wire N__41731;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41718;
    wire N__41711;
    wire N__41708;
    wire N__41707;
    wire N__41706;
    wire N__41705;
    wire N__41702;
    wire N__41699;
    wire N__41698;
    wire N__41693;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41674;
    wire N__41669;
    wire N__41666;
    wire N__41665;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41645;
    wire N__41644;
    wire N__41643;
    wire N__41642;
    wire N__41639;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41624;
    wire N__41619;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41603;
    wire N__41600;
    wire N__41599;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41579;
    wire N__41576;
    wire N__41575;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41555;
    wire N__41554;
    wire N__41551;
    wire N__41550;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41519;
    wire N__41516;
    wire N__41515;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41488;
    wire N__41487;
    wire N__41484;
    wire N__41479;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41467;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41447;
    wire N__41446;
    wire N__41443;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41420;
    wire N__41417;
    wire N__41416;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41396;
    wire N__41395;
    wire N__41392;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41362;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41352;
    wire N__41349;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41273;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41249;
    wire N__41248;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41231;
    wire N__41228;
    wire N__41227;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41207;
    wire N__41206;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41181;
    wire N__41174;
    wire N__41171;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41057;
    wire N__41054;
    wire N__41051;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41027;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41019;
    wire N__41014;
    wire N__41011;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40940;
    wire N__40937;
    wire N__40934;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40886;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40852;
    wire N__40851;
    wire N__40850;
    wire N__40849;
    wire N__40848;
    wire N__40847;
    wire N__40846;
    wire N__40845;
    wire N__40844;
    wire N__40843;
    wire N__40842;
    wire N__40839;
    wire N__40832;
    wire N__40831;
    wire N__40822;
    wire N__40817;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40795;
    wire N__40794;
    wire N__40793;
    wire N__40792;
    wire N__40791;
    wire N__40790;
    wire N__40789;
    wire N__40788;
    wire N__40787;
    wire N__40786;
    wire N__40785;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40762;
    wire N__40745;
    wire N__40730;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40724;
    wire N__40723;
    wire N__40722;
    wire N__40721;
    wire N__40720;
    wire N__40719;
    wire N__40718;
    wire N__40717;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40702;
    wire N__40701;
    wire N__40700;
    wire N__40699;
    wire N__40698;
    wire N__40697;
    wire N__40696;
    wire N__40695;
    wire N__40694;
    wire N__40693;
    wire N__40688;
    wire N__40685;
    wire N__40684;
    wire N__40683;
    wire N__40682;
    wire N__40681;
    wire N__40672;
    wire N__40671;
    wire N__40670;
    wire N__40667;
    wire N__40666;
    wire N__40659;
    wire N__40654;
    wire N__40653;
    wire N__40652;
    wire N__40649;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40615;
    wire N__40612;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40592;
    wire N__40587;
    wire N__40582;
    wire N__40577;
    wire N__40570;
    wire N__40559;
    wire N__40558;
    wire N__40555;
    wire N__40554;
    wire N__40553;
    wire N__40552;
    wire N__40551;
    wire N__40548;
    wire N__40547;
    wire N__40546;
    wire N__40541;
    wire N__40538;
    wire N__40537;
    wire N__40536;
    wire N__40535;
    wire N__40534;
    wire N__40533;
    wire N__40532;
    wire N__40531;
    wire N__40530;
    wire N__40529;
    wire N__40526;
    wire N__40525;
    wire N__40524;
    wire N__40521;
    wire N__40520;
    wire N__40519;
    wire N__40512;
    wire N__40511;
    wire N__40510;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40502;
    wire N__40499;
    wire N__40498;
    wire N__40497;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40489;
    wire N__40488;
    wire N__40487;
    wire N__40486;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40478;
    wire N__40477;
    wire N__40476;
    wire N__40475;
    wire N__40472;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40464;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40458;
    wire N__40445;
    wire N__40442;
    wire N__40437;
    wire N__40434;
    wire N__40429;
    wire N__40418;
    wire N__40407;
    wire N__40390;
    wire N__40385;
    wire N__40374;
    wire N__40371;
    wire N__40362;
    wire N__40359;
    wire N__40358;
    wire N__40355;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40318;
    wire N__40307;
    wire N__40304;
    wire N__40301;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40244;
    wire N__40243;
    wire N__40242;
    wire N__40241;
    wire N__40240;
    wire N__40239;
    wire N__40238;
    wire N__40237;
    wire N__40236;
    wire N__40235;
    wire N__40234;
    wire N__40233;
    wire N__40232;
    wire N__40231;
    wire N__40230;
    wire N__40229;
    wire N__40220;
    wire N__40203;
    wire N__40202;
    wire N__40201;
    wire N__40200;
    wire N__40199;
    wire N__40198;
    wire N__40197;
    wire N__40194;
    wire N__40193;
    wire N__40188;
    wire N__40185;
    wire N__40184;
    wire N__40179;
    wire N__40176;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40136;
    wire N__40127;
    wire N__40126;
    wire N__40125;
    wire N__40124;
    wire N__40123;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40117;
    wire N__40116;
    wire N__40115;
    wire N__40114;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40090;
    wire N__40087;
    wire N__40070;
    wire N__40067;
    wire N__40066;
    wire N__40065;
    wire N__40064;
    wire N__40063;
    wire N__40062;
    wire N__40061;
    wire N__40060;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40040;
    wire N__40029;
    wire N__40026;
    wire N__40025;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40006;
    wire N__40001;
    wire N__39996;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39964;
    wire N__39963;
    wire N__39962;
    wire N__39961;
    wire N__39960;
    wire N__39959;
    wire N__39958;
    wire N__39957;
    wire N__39956;
    wire N__39955;
    wire N__39954;
    wire N__39953;
    wire N__39952;
    wire N__39951;
    wire N__39950;
    wire N__39949;
    wire N__39948;
    wire N__39939;
    wire N__39938;
    wire N__39937;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39923;
    wire N__39920;
    wire N__39917;
    wire N__39916;
    wire N__39915;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39870;
    wire N__39865;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39847;
    wire N__39836;
    wire N__39833;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39818;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39784;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39759;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39740;
    wire N__39737;
    wire N__39728;
    wire N__39725;
    wire N__39724;
    wire N__39723;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39712;
    wire N__39709;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39690;
    wire N__39687;
    wire N__39682;
    wire N__39677;
    wire N__39674;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39659;
    wire N__39656;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39620;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39608;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39596;
    wire N__39593;
    wire N__39592;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39551;
    wire N__39550;
    wire N__39549;
    wire N__39548;
    wire N__39547;
    wire N__39546;
    wire N__39545;
    wire N__39544;
    wire N__39543;
    wire N__39542;
    wire N__39541;
    wire N__39540;
    wire N__39539;
    wire N__39538;
    wire N__39537;
    wire N__39536;
    wire N__39527;
    wire N__39518;
    wire N__39517;
    wire N__39516;
    wire N__39515;
    wire N__39514;
    wire N__39513;
    wire N__39512;
    wire N__39511;
    wire N__39510;
    wire N__39509;
    wire N__39508;
    wire N__39507;
    wire N__39506;
    wire N__39505;
    wire N__39504;
    wire N__39495;
    wire N__39486;
    wire N__39481;
    wire N__39472;
    wire N__39467;
    wire N__39458;
    wire N__39449;
    wire N__39444;
    wire N__39435;
    wire N__39428;
    wire N__39425;
    wire N__39424;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39406;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39353;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39337;
    wire N__39332;
    wire N__39329;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39221;
    wire N__39220;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39206;
    wire N__39205;
    wire N__39202;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39179;
    wire N__39176;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39128;
    wire N__39127;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39104;
    wire N__39103;
    wire N__39102;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39090;
    wire N__39087;
    wire N__39080;
    wire N__39077;
    wire N__39074;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38788;
    wire N__38785;
    wire N__38782;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38767;
    wire N__38764;
    wire N__38761;
    wire N__38758;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38698;
    wire N__38697;
    wire N__38692;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38682;
    wire N__38681;
    wire N__38680;
    wire N__38677;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38651;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38555;
    wire N__38552;
    wire N__38549;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38387;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38191;
    wire N__38190;
    wire N__38189;
    wire N__38186;
    wire N__38183;
    wire N__38180;
    wire N__38177;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38131;
    wire N__38130;
    wire N__38129;
    wire N__38126;
    wire N__38125;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38121;
    wire N__38120;
    wire N__38119;
    wire N__38118;
    wire N__38117;
    wire N__38116;
    wire N__38115;
    wire N__38114;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38106;
    wire N__38105;
    wire N__38104;
    wire N__38089;
    wire N__38072;
    wire N__38063;
    wire N__38062;
    wire N__38059;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38048;
    wire N__38047;
    wire N__38042;
    wire N__38039;
    wire N__38034;
    wire N__38031;
    wire N__38026;
    wire N__38015;
    wire N__38014;
    wire N__38013;
    wire N__38012;
    wire N__38011;
    wire N__38010;
    wire N__38009;
    wire N__38008;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37994;
    wire N__37993;
    wire N__37992;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37981;
    wire N__37980;
    wire N__37979;
    wire N__37978;
    wire N__37975;
    wire N__37974;
    wire N__37973;
    wire N__37972;
    wire N__37969;
    wire N__37952;
    wire N__37939;
    wire N__37938;
    wire N__37935;
    wire N__37934;
    wire N__37933;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37921;
    wire N__37914;
    wire N__37905;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37874;
    wire N__37873;
    wire N__37872;
    wire N__37871;
    wire N__37870;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37862;
    wire N__37861;
    wire N__37860;
    wire N__37859;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37845;
    wire N__37844;
    wire N__37843;
    wire N__37842;
    wire N__37841;
    wire N__37840;
    wire N__37839;
    wire N__37838;
    wire N__37833;
    wire N__37822;
    wire N__37813;
    wire N__37804;
    wire N__37799;
    wire N__37794;
    wire N__37793;
    wire N__37792;
    wire N__37791;
    wire N__37786;
    wire N__37781;
    wire N__37780;
    wire N__37775;
    wire N__37774;
    wire N__37769;
    wire N__37766;
    wire N__37761;
    wire N__37758;
    wire N__37755;
    wire N__37752;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37729;
    wire N__37726;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37649;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37321;
    wire N__37318;
    wire N__37315;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37030;
    wire N__37027;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37017;
    wire N__37010;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36953;
    wire N__36950;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36823;
    wire N__36820;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36805;
    wire N__36800;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36792;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36767;
    wire N__36764;
    wire N__36763;
    wire N__36762;
    wire N__36759;
    wire N__36754;
    wire N__36751;
    wire N__36746;
    wire N__36743;
    wire N__36742;
    wire N__36741;
    wire N__36738;
    wire N__36733;
    wire N__36728;
    wire N__36725;
    wire N__36724;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36709;
    wire N__36704;
    wire N__36701;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36693;
    wire N__36686;
    wire N__36681;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36650;
    wire N__36647;
    wire N__36646;
    wire N__36645;
    wire N__36642;
    wire N__36637;
    wire N__36634;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36598;
    wire N__36597;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36585;
    wire N__36582;
    wire N__36575;
    wire N__36574;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36536;
    wire N__36535;
    wire N__36534;
    wire N__36531;
    wire N__36526;
    wire N__36525;
    wire N__36520;
    wire N__36517;
    wire N__36512;
    wire N__36509;
    wire N__36508;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36491;
    wire N__36490;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36441;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36419;
    wire N__36418;
    wire N__36417;
    wire N__36414;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36374;
    wire N__36365;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36318;
    wire N__36317;
    wire N__36316;
    wire N__36315;
    wire N__36312;
    wire N__36295;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36291;
    wire N__36290;
    wire N__36289;
    wire N__36288;
    wire N__36287;
    wire N__36280;
    wire N__36279;
    wire N__36278;
    wire N__36273;
    wire N__36256;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36245;
    wire N__36240;
    wire N__36237;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36216;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36205;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36197;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36184;
    wire N__36183;
    wire N__36182;
    wire N__36181;
    wire N__36180;
    wire N__36177;
    wire N__36176;
    wire N__36173;
    wire N__36156;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36148;
    wire N__36145;
    wire N__36144;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36126;
    wire N__36109;
    wire N__36106;
    wire N__36105;
    wire N__36104;
    wire N__36103;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36091;
    wire N__36088;
    wire N__36081;
    wire N__36078;
    wire N__36065;
    wire N__36064;
    wire N__36063;
    wire N__36062;
    wire N__36061;
    wire N__36060;
    wire N__36057;
    wire N__36056;
    wire N__36055;
    wire N__36054;
    wire N__36053;
    wire N__36052;
    wire N__36051;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36036;
    wire N__36035;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36021;
    wire N__36018;
    wire N__36017;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36003;
    wire N__36002;
    wire N__36001;
    wire N__36000;
    wire N__35991;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35951;
    wire N__35942;
    wire N__35933;
    wire N__35930;
    wire N__35925;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35880;
    wire N__35879;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35841;
    wire N__35838;
    wire N__35837;
    wire N__35836;
    wire N__35833;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35813;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35617;
    wire N__35616;
    wire N__35615;
    wire N__35612;
    wire N__35611;
    wire N__35610;
    wire N__35605;
    wire N__35604;
    wire N__35601;
    wire N__35600;
    wire N__35599;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35587;
    wire N__35586;
    wire N__35585;
    wire N__35584;
    wire N__35583;
    wire N__35580;
    wire N__35577;
    wire N__35568;
    wire N__35559;
    wire N__35556;
    wire N__35547;
    wire N__35544;
    wire N__35543;
    wire N__35542;
    wire N__35541;
    wire N__35540;
    wire N__35537;
    wire N__35528;
    wire N__35525;
    wire N__35516;
    wire N__35513;
    wire N__35508;
    wire N__35501;
    wire N__35500;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35489;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35462;
    wire N__35453;
    wire N__35452;
    wire N__35451;
    wire N__35450;
    wire N__35449;
    wire N__35448;
    wire N__35447;
    wire N__35440;
    wire N__35439;
    wire N__35438;
    wire N__35437;
    wire N__35436;
    wire N__35427;
    wire N__35424;
    wire N__35415;
    wire N__35414;
    wire N__35413;
    wire N__35412;
    wire N__35409;
    wire N__35404;
    wire N__35397;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35368;
    wire N__35365;
    wire N__35364;
    wire N__35361;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35350;
    wire N__35347;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35315;
    wire N__35312;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35279;
    wire N__35278;
    wire N__35275;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35253;
    wire N__35252;
    wire N__35249;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35214;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35202;
    wire N__35195;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35180;
    wire N__35177;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35151;
    wire N__35144;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35136;
    wire N__35133;
    wire N__35132;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35105;
    wire N__35096;
    wire N__35095;
    wire N__35092;
    wire N__35091;
    wire N__35090;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35075;
    wire N__35072;
    wire N__35067;
    wire N__35064;
    wire N__35057;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35046;
    wire N__35045;
    wire N__35040;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35015;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35011;
    wire N__35010;
    wire N__35009;
    wire N__35002;
    wire N__34993;
    wire N__34992;
    wire N__34991;
    wire N__34990;
    wire N__34989;
    wire N__34988;
    wire N__34987;
    wire N__34986;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34969;
    wire N__34964;
    wire N__34963;
    wire N__34958;
    wire N__34955;
    wire N__34950;
    wire N__34949;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34925;
    wire N__34922;
    wire N__34915;
    wire N__34904;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34893;
    wire N__34888;
    wire N__34885;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34796;
    wire N__34793;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34775;
    wire N__34772;
    wire N__34771;
    wire N__34770;
    wire N__34769;
    wire N__34768;
    wire N__34765;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34742;
    wire N__34741;
    wire N__34738;
    wire N__34737;
    wire N__34736;
    wire N__34733;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34698;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34673;
    wire N__34672;
    wire N__34669;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34649;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34641;
    wire N__34640;
    wire N__34637;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34616;
    wire N__34607;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34596;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34565;
    wire N__34562;
    wire N__34561;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34543;
    wire N__34540;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34517;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34492;
    wire N__34487;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34451;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34439;
    wire N__34436;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34412;
    wire N__34411;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34379;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34371;
    wire N__34368;
    wire N__34363;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34345;
    wire N__34342;
    wire N__34341;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34329;
    wire N__34322;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34314;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34298;
    wire N__34295;
    wire N__34294;
    wire N__34293;
    wire N__34292;
    wire N__34287;
    wire N__34286;
    wire N__34285;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34252;
    wire N__34249;
    wire N__34248;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34227;
    wire N__34220;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34201;
    wire N__34196;
    wire N__34193;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34177;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34145;
    wire N__34142;
    wire N__34141;
    wire N__34140;
    wire N__34137;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34123;
    wire N__34120;
    wire N__34113;
    wire N__34110;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33950;
    wire N__33949;
    wire N__33946;
    wire N__33945;
    wire N__33942;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33930;
    wire N__33927;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33884;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33872;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33864;
    wire N__33861;
    wire N__33856;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33817;
    wire N__33814;
    wire N__33813;
    wire N__33806;
    wire N__33803;
    wire N__33802;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33778;
    wire N__33775;
    wire N__33774;
    wire N__33771;
    wire N__33766;
    wire N__33761;
    wire N__33760;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33731;
    wire N__33730;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33722;
    wire N__33719;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33688;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33565;
    wire N__33562;
    wire N__33561;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33504;
    wire N__33499;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33131;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33082;
    wire N__33081;
    wire N__33080;
    wire N__33079;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33073;
    wire N__33070;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33066;
    wire N__33065;
    wire N__33064;
    wire N__33063;
    wire N__33062;
    wire N__33045;
    wire N__33042;
    wire N__33041;
    wire N__33038;
    wire N__33037;
    wire N__33036;
    wire N__33035;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33015;
    wire N__33012;
    wire N__33011;
    wire N__33010;
    wire N__33009;
    wire N__33008;
    wire N__33007;
    wire N__33006;
    wire N__33005;
    wire N__33004;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32971;
    wire N__32968;
    wire N__32963;
    wire N__32958;
    wire N__32955;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32939;
    wire N__32926;
    wire N__32909;
    wire N__32908;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32892;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32881;
    wire N__32870;
    wire N__32865;
    wire N__32864;
    wire N__32863;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32859;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32841;
    wire N__32840;
    wire N__32839;
    wire N__32838;
    wire N__32837;
    wire N__32836;
    wire N__32835;
    wire N__32834;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32826;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32815;
    wire N__32812;
    wire N__32811;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32799;
    wire N__32790;
    wire N__32783;
    wire N__32770;
    wire N__32753;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32722;
    wire N__32721;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32711;
    wire N__32710;
    wire N__32709;
    wire N__32708;
    wire N__32707;
    wire N__32706;
    wire N__32705;
    wire N__32704;
    wire N__32703;
    wire N__32698;
    wire N__32695;
    wire N__32694;
    wire N__32693;
    wire N__32692;
    wire N__32691;
    wire N__32688;
    wire N__32671;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32648;
    wire N__32639;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32618;
    wire N__32613;
    wire N__32610;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32566;
    wire N__32561;
    wire N__32560;
    wire N__32559;
    wire N__32556;
    wire N__32555;
    wire N__32554;
    wire N__32553;
    wire N__32552;
    wire N__32551;
    wire N__32550;
    wire N__32549;
    wire N__32548;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32514;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32497;
    wire N__32492;
    wire N__32491;
    wire N__32490;
    wire N__32489;
    wire N__32486;
    wire N__32485;
    wire N__32484;
    wire N__32481;
    wire N__32480;
    wire N__32477;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32456;
    wire N__32453;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32404;
    wire N__32401;
    wire N__32396;
    wire N__32393;
    wire N__32384;
    wire N__32381;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32358;
    wire N__32349;
    wire N__32344;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32306;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32254;
    wire N__32249;
    wire N__32246;
    wire N__32245;
    wire N__32240;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32204;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32168;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32048;
    wire N__32047;
    wire N__32044;
    wire N__32041;
    wire N__32040;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32009;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31994;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31986;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31955;
    wire N__31954;
    wire N__31953;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31910;
    wire N__31907;
    wire N__31906;
    wire N__31901;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31865;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31829;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31719;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31683;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31654;
    wire N__31649;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31621;
    wire N__31616;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31591;
    wire N__31586;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31487;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31470;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31434;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31402;
    wire N__31397;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31382;
    wire N__31379;
    wire N__31376;
    wire N__31373;
    wire N__31372;
    wire N__31367;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31337;
    wire N__31336;
    wire N__31333;
    wire N__31332;
    wire N__31329;
    wire N__31324;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31275;
    wire N__31272;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31242;
    wire N__31235;
    wire N__31232;
    wire N__31231;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31220;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31193;
    wire N__31190;
    wire N__31189;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31145;
    wire N__31142;
    wire N__31141;
    wire N__31140;
    wire N__31137;
    wire N__31132;
    wire N__31129;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31018;
    wire N__31017;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30988;
    wire N__30987;
    wire N__30982;
    wire N__30979;
    wire N__30976;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30947;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30911;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30886;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30871;
    wire N__30868;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30850;
    wire N__30845;
    wire N__30844;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30827;
    wire N__30824;
    wire N__30819;
    wire N__30816;
    wire N__30809;
    wire N__30806;
    wire N__30805;
    wire N__30802;
    wire N__30801;
    wire N__30798;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30764;
    wire N__30763;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30746;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30697;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30661;
    wire N__30656;
    wire N__30655;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30624;
    wire N__30621;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30597;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30571;
    wire N__30566;
    wire N__30563;
    wire N__30562;
    wire N__30561;
    wire N__30556;
    wire N__30553;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30508;
    wire N__30507;
    wire N__30506;
    wire N__30503;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30470;
    wire N__30467;
    wire N__30466;
    wire N__30465;
    wire N__30460;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30403;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30349;
    wire N__30348;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30301;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30289;
    wire N__30286;
    wire N__30285;
    wire N__30282;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30248;
    wire N__30247;
    wire N__30246;
    wire N__30245;
    wire N__30244;
    wire N__30237;
    wire N__30234;
    wire N__30233;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30210;
    wire N__30203;
    wire N__30202;
    wire N__30199;
    wire N__30198;
    wire N__30195;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30164;
    wire N__30161;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30105;
    wire N__30104;
    wire N__30101;
    wire N__30096;
    wire N__30093;
    wire N__30086;
    wire N__30083;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30068;
    wire N__30065;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29948;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29764;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29694;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29659;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29633;
    wire N__29632;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29615;
    wire N__29612;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29538;
    wire N__29535;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29509;
    wire N__29508;
    wire N__29507;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29499;
    wire N__29496;
    wire N__29495;
    wire N__29492;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29423;
    wire N__29422;
    wire N__29419;
    wire N__29418;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29343;
    wire N__29336;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29296;
    wire N__29293;
    wire N__29292;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29258;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29218;
    wire N__29217;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29193;
    wire N__29186;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29079;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29046;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29024;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28984;
    wire N__28981;
    wire N__28980;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28955;
    wire N__28952;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28906;
    wire N__28903;
    wire N__28902;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28877;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28837;
    wire N__28834;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28793;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28747;
    wire N__28744;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28719;
    wire N__28712;
    wire N__28709;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28663;
    wire N__28660;
    wire N__28659;
    wire N__28656;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28634;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28591;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28563;
    wire N__28556;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28510;
    wire N__28509;
    wire N__28506;
    wire N__28505;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28484;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28441;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28424;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28412;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28366;
    wire N__28365;
    wire N__28362;
    wire N__28361;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28340;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28286;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28270;
    wire N__28265;
    wire N__28262;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28196;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28184;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28134;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28109;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28051;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28034;
    wire N__28031;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27965;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27922;
    wire N__27919;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27899;
    wire N__27896;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27809;
    wire N__27806;
    wire N__27805;
    wire N__27804;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27760;
    wire N__27755;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27691;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27568;
    wire N__27567;
    wire N__27564;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27518;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27507;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27473;
    wire N__27472;
    wire N__27471;
    wire N__27470;
    wire N__27467;
    wire N__27462;
    wire N__27459;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27447;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27358;
    wire N__27357;
    wire N__27356;
    wire N__27355;
    wire N__27354;
    wire N__27353;
    wire N__27352;
    wire N__27351;
    wire N__27350;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27342;
    wire N__27341;
    wire N__27340;
    wire N__27339;
    wire N__27338;
    wire N__27337;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27333;
    wire N__27332;
    wire N__27331;
    wire N__27330;
    wire N__27325;
    wire N__27316;
    wire N__27307;
    wire N__27298;
    wire N__27289;
    wire N__27280;
    wire N__27271;
    wire N__27262;
    wire N__27255;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27169;
    wire N__27164;
    wire N__27161;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27135;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27087;
    wire N__27082;
    wire N__27079;
    wire N__27068;
    wire N__27065;
    wire N__27064;
    wire N__27059;
    wire N__27056;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27044;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27038;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27011;
    wire N__27008;
    wire N__27007;
    wire N__27002;
    wire N__27001;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26952;
    wire N__26951;
    wire N__26948;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26914;
    wire N__26913;
    wire N__26912;
    wire N__26909;
    wire N__26904;
    wire N__26901;
    wire N__26896;
    wire N__26893;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26874;
    wire N__26869;
    wire N__26868;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26840;
    wire N__26837;
    wire N__26832;
    wire N__26829;
    wire N__26824;
    wire N__26821;
    wire N__26816;
    wire N__26813;
    wire N__26812;
    wire N__26807;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26799;
    wire N__26794;
    wire N__26791;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26770;
    wire N__26769;
    wire N__26766;
    wire N__26765;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26738;
    wire N__26735;
    wire N__26734;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26720;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26704;
    wire N__26701;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26681;
    wire N__26678;
    wire N__26673;
    wire N__26670;
    wire N__26665;
    wire N__26662;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26644;
    wire N__26643;
    wire N__26640;
    wire N__26635;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26599;
    wire N__26598;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26578;
    wire N__26575;
    wire N__26570;
    wire N__26567;
    wire N__26566;
    wire N__26565;
    wire N__26562;
    wire N__26557;
    wire N__26556;
    wire N__26551;
    wire N__26548;
    wire N__26543;
    wire N__26540;
    wire N__26539;
    wire N__26538;
    wire N__26535;
    wire N__26530;
    wire N__26525;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26489;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26459;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26402;
    wire N__26399;
    wire N__26398;
    wire N__26397;
    wire N__26394;
    wire N__26389;
    wire N__26388;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26368;
    wire N__26367;
    wire N__26366;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26320;
    wire N__26317;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26305;
    wire N__26304;
    wire N__26303;
    wire N__26300;
    wire N__26295;
    wire N__26292;
    wire N__26287;
    wire N__26284;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26232;
    wire N__26229;
    wire N__26224;
    wire N__26219;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26194;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26161;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26146;
    wire N__26141;
    wire N__26140;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26113;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26101;
    wire N__26098;
    wire N__26097;
    wire N__26090;
    wire N__26087;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26069;
    wire N__26068;
    wire N__26067;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26049;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26023;
    wire N__26020;
    wire N__26019;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25994;
    wire N__25991;
    wire N__25990;
    wire N__25989;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25933;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25918;
    wire N__25915;
    wire N__25910;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25891;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25880;
    wire N__25877;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25837;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25826;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25798;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25770;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25754;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25739;
    wire N__25736;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25711;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25681;
    wire N__25680;
    wire N__25677;
    wire N__25676;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25657;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25642;
    wire N__25641;
    wire N__25634;
    wire N__25631;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25613;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25605;
    wire N__25602;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25573;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25504;
    wire N__25503;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25488;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25264;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24967;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24928;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24908;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24900;
    wire N__24897;
    wire N__24892;
    wire N__24887;
    wire N__24884;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24490;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24409;
    wire N__24406;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24389;
    wire N__24388;
    wire N__24385;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24368;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24344;
    wire N__24341;
    wire N__24340;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24299;
    wire N__24298;
    wire N__24297;
    wire N__24296;
    wire N__24295;
    wire N__24294;
    wire N__24293;
    wire N__24292;
    wire N__24291;
    wire N__24290;
    wire N__24281;
    wire N__24272;
    wire N__24267;
    wire N__24262;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24236;
    wire N__24235;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24218;
    wire N__24217;
    wire N__24214;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24116;
    wire N__24113;
    wire N__24112;
    wire N__24109;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24094;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24082;
    wire N__24081;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24034;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__24001;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23986;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23966;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23961;
    wire N__23960;
    wire N__23959;
    wire N__23958;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23954;
    wire N__23953;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23947;
    wire N__23946;
    wire N__23945;
    wire N__23944;
    wire N__23943;
    wire N__23942;
    wire N__23941;
    wire N__23940;
    wire N__23931;
    wire N__23922;
    wire N__23913;
    wire N__23904;
    wire N__23895;
    wire N__23886;
    wire N__23881;
    wire N__23872;
    wire N__23867;
    wire N__23858;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23812;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23779;
    wire N__23774;
    wire N__23771;
    wire N__23770;
    wire N__23769;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23735;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23720;
    wire N__23717;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23690;
    wire N__23687;
    wire N__23686;
    wire N__23681;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23666;
    wire N__23663;
    wire N__23662;
    wire N__23661;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23638;
    wire N__23635;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23620;
    wire N__23615;
    wire N__23612;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23579;
    wire N__23576;
    wire N__23575;
    wire N__23572;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23557;
    wire N__23552;
    wire N__23549;
    wire N__23548;
    wire N__23547;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23520;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23504;
    wire N__23501;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23489;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23460;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23444;
    wire N__23441;
    wire N__23440;
    wire N__23435;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23420;
    wire N__23417;
    wire N__23416;
    wire N__23415;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23392;
    wire N__23389;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23374;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23355;
    wire N__23350;
    wire N__23347;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23328;
    wire N__23323;
    wire N__23320;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23308;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23293;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23274;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23258;
    wire N__23255;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23243;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23228;
    wire N__23225;
    wire N__23224;
    wire N__23219;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23204;
    wire N__23201;
    wire N__23200;
    wire N__23195;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23180;
    wire N__23177;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23162;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23122;
    wire N__23121;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23094;
    wire N__23093;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23085;
    wire N__23084;
    wire N__23081;
    wire N__23074;
    wire N__23065;
    wire N__23064;
    wire N__23063;
    wire N__23062;
    wire N__23061;
    wire N__23060;
    wire N__23059;
    wire N__23058;
    wire N__23057;
    wire N__23056;
    wire N__23055;
    wire N__23052;
    wire N__23051;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23036;
    wire N__23035;
    wire N__23034;
    wire N__23033;
    wire N__23032;
    wire N__23031;
    wire N__23030;
    wire N__23029;
    wire N__23028;
    wire N__23027;
    wire N__23020;
    wire N__23017;
    wire N__23010;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22982;
    wire N__22975;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22921;
    wire N__22918;
    wire N__22913;
    wire N__22906;
    wire N__22897;
    wire N__22890;
    wire N__22879;
    wire N__22878;
    wire N__22877;
    wire N__22876;
    wire N__22875;
    wire N__22874;
    wire N__22863;
    wire N__22860;
    wire N__22859;
    wire N__22858;
    wire N__22857;
    wire N__22854;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22809;
    wire N__22804;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22781;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22754;
    wire N__22749;
    wire N__22742;
    wire N__22741;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22723;
    wire N__22720;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22639;
    wire N__22636;
    wire N__22635;
    wire N__22634;
    wire N__22631;
    wire N__22626;
    wire N__22623;
    wire N__22616;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22608;
    wire N__22603;
    wire N__22600;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22387;
    wire N__22386;
    wire N__22385;
    wire N__22384;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22150;
    wire N__22149;
    wire N__22148;
    wire N__22147;
    wire N__22144;
    wire N__22143;
    wire N__22140;
    wire N__22139;
    wire N__22136;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22096;
    wire N__22093;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22071;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21862;
    wire N__21861;
    wire N__21860;
    wire N__21855;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21825;
    wire N__21818;
    wire N__21815;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21704;
    wire N__21701;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21686;
    wire N__21683;
    wire N__21682;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21643;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21574;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21556;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21514;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21493;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21452;
    wire N__21449;
    wire N__21448;
    wire N__21445;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21410;
    wire N__21407;
    wire N__21406;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21349;
    wire N__21344;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21310;
    wire N__21307;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21279;
    wire N__21274;
    wire N__21271;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21212;
    wire N__21209;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21160;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21106;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21091;
    wire N__21090;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21084;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21059;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21051;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21026;
    wire N__21025;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21005;
    wire N__20998;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20885;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20859;
    wire N__20854;
    wire N__20851;
    wire N__20846;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20792;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20780;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20705;
    wire N__20704;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20678;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20615;
    wire N__20614;
    wire N__20613;
    wire N__20612;
    wire N__20611;
    wire N__20610;
    wire N__20609;
    wire N__20608;
    wire N__20607;
    wire N__20606;
    wire N__20605;
    wire N__20604;
    wire N__20603;
    wire N__20602;
    wire N__20601;
    wire N__20600;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20574;
    wire N__20559;
    wire N__20558;
    wire N__20557;
    wire N__20556;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20548;
    wire N__20545;
    wire N__20540;
    wire N__20537;
    wire N__20532;
    wire N__20531;
    wire N__20530;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20503;
    wire N__20500;
    wire N__20493;
    wire N__20488;
    wire N__20483;
    wire N__20474;
    wire N__20471;
    wire N__20466;
    wire N__20463;
    wire N__20450;
    wire N__20449;
    wire N__20448;
    wire N__20447;
    wire N__20446;
    wire N__20445;
    wire N__20432;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20422;
    wire N__20421;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20409;
    wire N__20402;
    wire N__20401;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20397;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20379;
    wire N__20378;
    wire N__20375;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20349;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20297;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20270;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20167;
    wire N__20164;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20098;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20037;
    wire N__20036;
    wire N__20035;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20031;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20012;
    wire N__20007;
    wire N__20004;
    wire N__19997;
    wire N__19996;
    wire N__19995;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19979;
    wire N__19974;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19891;
    wire N__19890;
    wire N__19889;
    wire N__19888;
    wire N__19887;
    wire N__19886;
    wire N__19885;
    wire N__19882;
    wire N__19877;
    wire N__19872;
    wire N__19867;
    wire N__19864;
    wire N__19863;
    wire N__19858;
    wire N__19855;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19839;
    wire N__19836;
    wire N__19829;
    wire N__19828;
    wire N__19827;
    wire N__19826;
    wire N__19823;
    wire N__19816;
    wire N__19815;
    wire N__19814;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19802;
    wire N__19799;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19780;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19675;
    wire N__19674;
    wire N__19673;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19665;
    wire N__19662;
    wire N__19661;
    wire N__19658;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19638;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19576;
    wire N__19575;
    wire N__19572;
    wire N__19567;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19504;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19015;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18986;
    wire N__18985;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18953;
    wire N__18952;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18909;
    wire N__18906;
    wire N__18901;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18868;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18839;
    wire N__18838;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18794;
    wire N__18791;
    wire N__18790;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18771;
    wire N__18766;
    wire N__18763;
    wire N__18758;
    wire N__18757;
    wire N__18756;
    wire N__18753;
    wire N__18748;
    wire N__18745;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18732;
    wire N__18729;
    wire N__18724;
    wire N__18721;
    wire N__18716;
    wire N__18713;
    wire N__18712;
    wire N__18711;
    wire N__18708;
    wire N__18703;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18691;
    wire N__18690;
    wire N__18687;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18668;
    wire N__18667;
    wire N__18666;
    wire N__18659;
    wire N__18656;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18644;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18632;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18349;
    wire N__18344;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18338;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_1_7_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_1_8_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire bfn_1_12_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire un7_start_stop_0_a3;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire pwm_duty_input_8;
    wire pwm_duty_input_9;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_2;
    wire pwm_duty_input_1;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire bfn_2_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_2_13_0_;
    wire N_32_i_i;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire bfn_3_8_0_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_178 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire bfn_4_5_0_;
    wire un5_counter_cry_1;
    wire un5_counter_cry_2;
    wire un5_counter_cry_3;
    wire un5_counter_cry_4;
    wire un5_counter_cry_5;
    wire un5_counter_cry_6;
    wire un5_counter_cry_7;
    wire un5_counter_cry_8;
    wire bfn_4_6_0_;
    wire un5_counter_cry_9;
    wire un5_counter_cry_10;
    wire un5_counter_cry_11;
    wire counterZ0Z_11;
    wire counterZ0Z_9;
    wire counterZ0Z_8;
    wire counterZ0Z_2;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire counter_RNO_0Z0Z_7;
    wire counterZ0Z_7;
    wire N_19_1;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire counterZ0Z_4;
    wire counterZ0Z_3;
    wire counterZ0Z_5;
    wire counterZ0Z_6;
    wire un2_counter_5_cascade_;
    wire counter_RNO_0Z0Z_12;
    wire counterZ0Z_12;
    wire counter_RNO_0Z0Z_10;
    wire counterZ0Z_10;
    wire counterZ0Z_1;
    wire counterZ0Z_0;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire un2_counter_8;
    wire un2_counter_7;
    wire un2_counter_9;
    wire clk_10khz_RNIIENAZ0Z2_cascade_;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_5_9_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_5_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_5_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_5_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire clk_10khz_i;
    wire clk_10khz_RNIIENAZ0Z2;
    wire \delay_measurement_inst.delay_hc_reg3lt19_0 ;
    wire \delay_measurement_inst.delay_hc_reg3lt19_0_cascade_ ;
    wire bfn_7_19_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ;
    wire bfn_7_20_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ;
    wire bfn_7_21_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ;
    wire bfn_7_22_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_phase.N_188_i_g ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_8_8_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_8_9_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_reg3lto31_5_0 ;
    wire bfn_8_13_0_;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire bfn_8_14_0_;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_input_1_cry_11 ;
    wire \current_shift_inst.control_input_1_cry_12 ;
    wire \current_shift_inst.control_input_1_cry_13 ;
    wire \current_shift_inst.control_input_1_cry_14 ;
    wire \current_shift_inst.control_input_1_cry_15 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.control_input_1_cry_16 ;
    wire \current_shift_inst.control_input_1_cry_17 ;
    wire \current_shift_inst.control_input_1_cry_18 ;
    wire \current_shift_inst.control_input_1_cry_19 ;
    wire \current_shift_inst.control_input_1_cry_20 ;
    wire \current_shift_inst.control_input_1_cry_21 ;
    wire \current_shift_inst.control_input_1_cry_22 ;
    wire \current_shift_inst.control_input_1_cry_23 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.control_input_1_cry_24 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_2 ;
    wire \current_shift_inst.z_5_cry_1 ;
    wire \current_shift_inst.elapsed_time_ns_phase_3 ;
    wire \current_shift_inst.z_5_cry_2 ;
    wire \current_shift_inst.z_5_cry_3 ;
    wire \current_shift_inst.z_5_cry_4 ;
    wire \current_shift_inst.z_5_cry_5 ;
    wire \current_shift_inst.z_5_cry_6 ;
    wire \current_shift_inst.z_5_cry_7 ;
    wire \current_shift_inst.z_5_cry_8 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.z_5_cry_9 ;
    wire \current_shift_inst.z_5_cry_10 ;
    wire \current_shift_inst.z_5_cry_11 ;
    wire \current_shift_inst.z_5_cry_12 ;
    wire \current_shift_inst.z_5_cry_13 ;
    wire \current_shift_inst.z_5_cry_14 ;
    wire \current_shift_inst.z_5_cry_15 ;
    wire \current_shift_inst.z_5_cry_16 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.z_5_cry_17 ;
    wire \current_shift_inst.z_5_cry_18 ;
    wire \current_shift_inst.z_5_cry_19 ;
    wire \current_shift_inst.z_5_cry_20 ;
    wire \current_shift_inst.z_5_cry_21 ;
    wire \current_shift_inst.z_5_cry_22 ;
    wire \current_shift_inst.z_5_cry_23 ;
    wire \current_shift_inst.z_5_cry_24 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.z_5_cry_25 ;
    wire \current_shift_inst.z_5_cry_26 ;
    wire \current_shift_inst.z_5_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_phase_29 ;
    wire \current_shift_inst.z_5_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.elapsed_time_ns_phase_30 ;
    wire \current_shift_inst.z_5_cry_29 ;
    wire \current_shift_inst.z_5_cry_30 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_0 ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_1 ;
    wire \current_shift_inst.timer_phase.counter_cry_0 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_2 ;
    wire \current_shift_inst.timer_phase.counter_cry_1 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_3 ;
    wire \current_shift_inst.timer_phase.counter_cry_2 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_4 ;
    wire \current_shift_inst.timer_phase.counter_cry_3 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_5 ;
    wire \current_shift_inst.timer_phase.counter_cry_4 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_6 ;
    wire \current_shift_inst.timer_phase.counter_cry_5 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_7 ;
    wire \current_shift_inst.timer_phase.counter_cry_6 ;
    wire \current_shift_inst.timer_phase.counter_cry_7 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_8 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_9 ;
    wire \current_shift_inst.timer_phase.counter_cry_8 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_10 ;
    wire \current_shift_inst.timer_phase.counter_cry_9 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_11 ;
    wire \current_shift_inst.timer_phase.counter_cry_10 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_12 ;
    wire \current_shift_inst.timer_phase.counter_cry_11 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_13 ;
    wire \current_shift_inst.timer_phase.counter_cry_12 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_14 ;
    wire \current_shift_inst.timer_phase.counter_cry_13 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_15 ;
    wire \current_shift_inst.timer_phase.counter_cry_14 ;
    wire \current_shift_inst.timer_phase.counter_cry_15 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_16 ;
    wire bfn_8_23_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_17 ;
    wire \current_shift_inst.timer_phase.counter_cry_16 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_18 ;
    wire \current_shift_inst.timer_phase.counter_cry_17 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_19 ;
    wire \current_shift_inst.timer_phase.counter_cry_18 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_20 ;
    wire \current_shift_inst.timer_phase.counter_cry_19 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_21 ;
    wire \current_shift_inst.timer_phase.counter_cry_20 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_22 ;
    wire \current_shift_inst.timer_phase.counter_cry_21 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_23 ;
    wire \current_shift_inst.timer_phase.counter_cry_22 ;
    wire \current_shift_inst.timer_phase.counter_cry_23 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_24 ;
    wire bfn_8_24_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_25 ;
    wire \current_shift_inst.timer_phase.counter_cry_24 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_26 ;
    wire \current_shift_inst.timer_phase.counter_cry_25 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_27 ;
    wire \current_shift_inst.timer_phase.counter_cry_26 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_28 ;
    wire \current_shift_inst.timer_phase.counter_cry_27 ;
    wire \current_shift_inst.timer_phase.counter_cry_28 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_187_i ;
    wire \current_shift_inst.timer_phase.N_193_i ;
    wire \current_shift_inst.timer_phase.running_i ;
    wire il_max_comp1_c;
    wire bfn_9_7_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_9_8_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.un1_counterlto2_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire bfn_9_13_0_;
    wire \current_shift_inst.z_i_0_31 ;
    wire \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ;
    wire \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_1 ;
    wire \current_shift_inst.N_1620_i ;
    wire \current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_4 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_6 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire bfn_9_14_0_;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_7 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_8 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_cry_9 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_10 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_0_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_cry_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_14 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.un38_control_input_0_cry_15 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_cry_16 ;
    wire \current_shift_inst.control_input_1_axb_12 ;
    wire \current_shift_inst.un38_control_input_0_cry_17 ;
    wire \current_shift_inst.control_input_1_axb_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_18 ;
    wire \current_shift_inst.control_input_1_axb_14 ;
    wire \current_shift_inst.un38_control_input_0_cry_19 ;
    wire \current_shift_inst.control_input_1_axb_15 ;
    wire \current_shift_inst.un38_control_input_0_cry_20 ;
    wire \current_shift_inst.control_input_1_axb_16 ;
    wire \current_shift_inst.un38_control_input_0_cry_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_22 ;
    wire \current_shift_inst.control_input_1_axb_17 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ;
    wire \current_shift_inst.control_input_1_axb_18 ;
    wire \current_shift_inst.un38_control_input_0_cry_23 ;
    wire \current_shift_inst.control_input_1_axb_19 ;
    wire \current_shift_inst.un38_control_input_0_cry_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ;
    wire \current_shift_inst.control_input_1_axb_20 ;
    wire \current_shift_inst.un38_control_input_0_cry_25 ;
    wire \current_shift_inst.control_input_1_axb_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ;
    wire \current_shift_inst.control_input_1_axb_22 ;
    wire \current_shift_inst.un38_control_input_0_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ;
    wire \current_shift_inst.control_input_1_axb_23 ;
    wire \current_shift_inst.un38_control_input_0_cry_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ;
    wire \current_shift_inst.control_input_1_axb_24 ;
    wire \current_shift_inst.un38_control_input_0_cry_29 ;
    wire \current_shift_inst.un38_control_input_0_cry_30 ;
    wire \current_shift_inst.un38_control_input_0_axb_31 ;
    wire \current_shift_inst.control_input_1_cry_24_THRU_CO ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.phase_valid_RNISLORZ0Z2 ;
    wire G_406;
    wire bfn_9_18_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_1 ;
    wire G_405;
    wire \current_shift_inst.z_cry_0 ;
    wire \current_shift_inst.z_5_2 ;
    wire \current_shift_inst.z_cry_1 ;
    wire \current_shift_inst.z_5_3 ;
    wire \current_shift_inst.z_cry_2 ;
    wire \current_shift_inst.z_5_4 ;
    wire \current_shift_inst.z_cry_3 ;
    wire \current_shift_inst.z_5_5 ;
    wire \current_shift_inst.z_cry_4 ;
    wire \current_shift_inst.z_5_6 ;
    wire \current_shift_inst.z_cry_5 ;
    wire \current_shift_inst.z_5_7 ;
    wire \current_shift_inst.z_cry_6 ;
    wire \current_shift_inst.z_cry_7 ;
    wire \current_shift_inst.z_5_8 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.z_5_9 ;
    wire \current_shift_inst.z_cry_8 ;
    wire \current_shift_inst.z_5_10 ;
    wire \current_shift_inst.z_cry_9 ;
    wire \current_shift_inst.z_5_11 ;
    wire \current_shift_inst.z_cry_10 ;
    wire \current_shift_inst.z_5_12 ;
    wire \current_shift_inst.z_cry_11 ;
    wire \current_shift_inst.z_5_13 ;
    wire \current_shift_inst.z_cry_12 ;
    wire \current_shift_inst.z_5_14 ;
    wire \current_shift_inst.z_cry_13 ;
    wire \current_shift_inst.z_5_15 ;
    wire \current_shift_inst.z_cry_14 ;
    wire \current_shift_inst.z_cry_15 ;
    wire \current_shift_inst.z_5_16 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.z_5_17 ;
    wire \current_shift_inst.z_cry_16 ;
    wire \current_shift_inst.z_5_18 ;
    wire \current_shift_inst.z_cry_17 ;
    wire \current_shift_inst.z_5_19 ;
    wire \current_shift_inst.z_cry_18 ;
    wire \current_shift_inst.z_5_20 ;
    wire \current_shift_inst.z_cry_19 ;
    wire \current_shift_inst.z_5_21 ;
    wire \current_shift_inst.z_cry_20 ;
    wire \current_shift_inst.z_5_22 ;
    wire \current_shift_inst.z_cry_21 ;
    wire \current_shift_inst.z_5_23 ;
    wire \current_shift_inst.z_cry_22 ;
    wire \current_shift_inst.z_cry_23 ;
    wire \current_shift_inst.z_5_24 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.z_5_25 ;
    wire \current_shift_inst.z_cry_24 ;
    wire \current_shift_inst.z_5_26 ;
    wire \current_shift_inst.z_cry_25 ;
    wire \current_shift_inst.z_5_27 ;
    wire \current_shift_inst.z_cry_26 ;
    wire \current_shift_inst.z_5_28 ;
    wire \current_shift_inst.z_cry_27 ;
    wire \current_shift_inst.z_5_29 ;
    wire \current_shift_inst.z_cry_28 ;
    wire \current_shift_inst.z_5_30 ;
    wire \current_shift_inst.z_cry_29 ;
    wire \current_shift_inst.z_5_cry_30_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_phase_31 ;
    wire \current_shift_inst.z_cry_30 ;
    wire \current_shift_inst.stop_timer_s1_RNOZ0Z_0 ;
    wire \current_shift_inst.start_timer_phaseZ0 ;
    wire il_max_comp1_D1;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILORI_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ;
    wire \current_shift_inst.elapsed_time_ns_phase_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ;
    wire \current_shift_inst.elapsed_time_ns_phase_5 ;
    wire \current_shift_inst.elapsed_time_ns_phase_4 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ;
    wire \current_shift_inst.elapsed_time_ns_phase_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ;
    wire \current_shift_inst.elapsed_time_ns_phase_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ;
    wire \current_shift_inst.elapsed_time_ns_phase_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ;
    wire \current_shift_inst.elapsed_time_ns_phase_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ;
    wire \current_shift_inst.elapsed_time_ns_phase_9 ;
    wire \current_shift_inst.elapsed_time_ns_phase_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ;
    wire \current_shift_inst.elapsed_time_ns_phase_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ;
    wire \current_shift_inst.elapsed_time_ns_phase_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ;
    wire \current_shift_inst.elapsed_time_ns_phase_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI190J_15 ;
    wire \current_shift_inst.elapsed_time_ns_phase_20 ;
    wire \current_shift_inst.elapsed_time_ns_phase_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ;
    wire \current_shift_inst.elapsed_time_ns_phase_17 ;
    wire \current_shift_inst.elapsed_time_ns_phase_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ;
    wire \current_shift_inst.un38_control_input_0 ;
    wire bfn_10_17_0_;
    wire \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_1 ;
    wire \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_2 ;
    wire \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_3 ;
    wire \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_4 ;
    wire \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_5 ;
    wire \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_6 ;
    wire \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_7 ;
    wire \current_shift_inst.un4_control_input_cry_8 ;
    wire \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ;
    wire bfn_10_18_0_;
    wire \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ;
    wire \current_shift_inst.un4_control_input_cry_9 ;
    wire \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_10 ;
    wire \current_shift_inst.un4_control_input_cry_11 ;
    wire \current_shift_inst.un4_control_input_cry_12 ;
    wire \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_13 ;
    wire \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_14 ;
    wire \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_15 ;
    wire \current_shift_inst.un4_control_input_cry_16 ;
    wire \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ;
    wire bfn_10_19_0_;
    wire \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_17 ;
    wire \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_18 ;
    wire \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_19 ;
    wire \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_20 ;
    wire \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_21 ;
    wire \current_shift_inst.un4_control_input_cry_22 ;
    wire \current_shift_inst.un4_control_input_cry_23 ;
    wire \current_shift_inst.un4_control_input_cry_24 ;
    wire bfn_10_20_0_;
    wire \current_shift_inst.un4_control_input_cry_25 ;
    wire \current_shift_inst.un4_control_input_cry_26 ;
    wire \current_shift_inst.un4_control_input_cry_27 ;
    wire \current_shift_inst.un4_control_input_cry_28 ;
    wire \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ;
    wire \current_shift_inst.un4_control_input_cry_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input_cry_30 ;
    wire \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_28 ;
    wire \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ;
    wire bfn_10_21_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire bfn_10_22_0_;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire bfn_10_23_0_;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire bfn_10_24_0_;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_192_i ;
    wire \current_shift_inst.timer_phase.runningZ0 ;
    wire \current_shift_inst.stop_timer_phaseZ0 ;
    wire \current_shift_inst.timer_phase.N_188_i ;
    wire il_max_comp2_c;
    wire il_min_comp2_c;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_axb_0 ;
    wire bfn_11_10_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire bfn_11_11_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.control_inputZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.control_inputZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.control_inputZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.control_inputZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.control_inputZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire bfn_11_12_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.control_inputZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.control_inputZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.control_inputZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.control_inputZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.control_inputZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.control_inputZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.control_inputZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.control_inputZ0Z_24 ;
    wire bfn_11_13_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.control_inputZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_fast_31 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input_axb_1 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input_axb_2 ;
    wire \current_shift_inst.un4_control_input_axb_14 ;
    wire \current_shift_inst.un4_control_input_axb_3 ;
    wire \current_shift_inst.un4_control_input_axb_4 ;
    wire \current_shift_inst.un4_control_input_axb_5 ;
    wire \current_shift_inst.un4_control_input_axb_6 ;
    wire \current_shift_inst.un4_control_input_axb_7 ;
    wire \current_shift_inst.un4_control_input_axb_8 ;
    wire \current_shift_inst.un4_control_input_axb_13 ;
    wire \current_shift_inst.un4_control_input_axb_15 ;
    wire \current_shift_inst.un4_control_input_axb_9 ;
    wire \current_shift_inst.un4_control_input_axb_10 ;
    wire \current_shift_inst.un4_control_input_axb_11 ;
    wire \current_shift_inst.un4_control_input_axb_12 ;
    wire \current_shift_inst.un4_control_input_axb_16 ;
    wire \current_shift_inst.un4_control_input_axb_20 ;
    wire \current_shift_inst.un4_control_input_axb_18 ;
    wire \current_shift_inst.un4_control_input_axb_23 ;
    wire \current_shift_inst.un4_control_input_axb_19 ;
    wire \current_shift_inst.un4_control_input_axb_25 ;
    wire \current_shift_inst.un4_control_input_axb_22 ;
    wire \current_shift_inst.un4_control_input_axb_24 ;
    wire \current_shift_inst.un4_control_input_axb_17 ;
    wire \current_shift_inst.un4_control_input_axb_21 ;
    wire \current_shift_inst.un4_control_input_axb_26 ;
    wire \current_shift_inst.z_31 ;
    wire \current_shift_inst.z_i_31 ;
    wire \current_shift_inst.un4_control_input_axb_30 ;
    wire \current_shift_inst.un4_control_input_axb_27 ;
    wire \current_shift_inst.un4_control_input_axb_29 ;
    wire \current_shift_inst.un4_control_input_axb_28 ;
    wire \current_shift_inst.S1_sync_prevZ0 ;
    wire \current_shift_inst.S1_syncZ0Z0 ;
    wire \current_shift_inst.S1_syncZ0Z1 ;
    wire \current_shift_inst.meas_stateZ0Z_0 ;
    wire \current_shift_inst.S1_riseZ0 ;
    wire \current_shift_inst.phase_validZ0 ;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire il_min_comp2_D1;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_20 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_m5_iZ0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_N_4_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_phase_11 ;
    wire \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ;
    wire \current_shift_inst.elapsed_time_ns_phase_27 ;
    wire \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ;
    wire \current_shift_inst.elapsed_time_ns_phase_23 ;
    wire \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ;
    wire \current_shift_inst.elapsed_time_ns_phase_22 ;
    wire \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ;
    wire \current_shift_inst.elapsed_time_ns_phase_26 ;
    wire \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ;
    wire \current_shift_inst.elapsed_time_ns_phase_24 ;
    wire \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ;
    wire bfn_12_19_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ;
    wire bfn_12_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ;
    wire bfn_12_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ;
    wire bfn_12_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_187_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire s1_phy_c;
    wire \current_shift_inst.S3_riseZ0 ;
    wire \current_shift_inst.S3_sync_prevZ0 ;
    wire \current_shift_inst.S3_syncZ0Z0 ;
    wire \current_shift_inst.S3_syncZ0Z1 ;
    wire il_max_comp2_D1;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.N_79 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire N_605_g;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_13_13_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_13_14_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_13_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire \phase_controller_slave.state_RNIVDE2Z0Z_0_cascade_ ;
    wire state_ns_i_a2_1;
    wire start_stop_c;
    wire s4_phy_c;
    wire il_min_comp2_D2;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_slave.state_RNIVDE2Z0Z_0 ;
    wire s3_phy_c;
    wire shift_flag_start;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire bfn_13_24_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_13_25_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_13_26_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire s2_phy_c;
    wire \delay_measurement_inst.delay_hc_timer.N_335_i ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ;
    wire measured_delay_hc_23;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_N_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0_cascade_ ;
    wire measured_delay_hc_16;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0 ;
    wire measured_delay_hc_17;
    wire measured_delay_hc_10;
    wire measured_delay_hc_11;
    wire measured_delay_hc_2;
    wire measured_delay_hc_7;
    wire measured_delay_hc_5;
    wire measured_delay_hc_12;
    wire measured_delay_hc_1;
    wire measured_delay_hc_3;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ;
    wire measured_delay_hc_15;
    wire measured_delay_hc_13;
    wire measured_delay_hc_18;
    wire measured_delay_hc_6;
    wire \phase_controller_inst1.stoper_hc.un1_startlt31_0 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31 ;
    wire measured_delay_hc_8;
    wire \phase_controller_inst1.stoper_hc.un1_start ;
    wire bfn_14_18_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_14_19_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_14_20_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire red_c_i;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire delay_tr_d2;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire delay_hc_d2;
    wire measured_delay_hc_9;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_ ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_c_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_0_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9 ;
    wire measured_delay_hc_21;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ;
    wire measured_delay_hc_20;
    wire measured_delay_hc_19;
    wire measured_delay_hc_22;
    wire \delay_measurement_inst.delay_hc_reg3lto31_0_0 ;
    wire measured_delay_hc_29;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ;
    wire measured_delay_hc_27;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_15_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire bfn_15_14_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_15_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_15_16_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire bfn_15_17_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire bfn_15_18_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_slave.stoper_tr.time_passed11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_21_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_22_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_15_23_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_24_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_25_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_15_26_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire bfn_16_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_16_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_16_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_16_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.N_336_i ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_reg3lto30_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_0 ;
    wire \delay_measurement_inst.delay_hc_reg3lto30_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_reg3_cascade_ ;
    wire measured_delay_hc_4;
    wire measured_delay_hc_14;
    wire measured_delay_hc_24;
    wire measured_delay_hc_25;
    wire measured_delay_hc_26;
    wire measured_delay_hc_28;
    wire measured_delay_hc_30;
    wire measured_delay_hc_0;
    wire \delay_measurement_inst.delay_hc_reg3 ;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire measured_delay_hc_31;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire measured_delay_tr_10;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire measured_delay_tr_12;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_17_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_17_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4Z0Z_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_7_0 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_17_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_17_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_17_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_338_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_293 ;
    wire \delay_measurement_inst.N_358_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ;
    wire \delay_measurement_inst.N_307 ;
    wire \phase_controller_slave.start_timer_hc_RNO_0_0 ;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_ ;
    wire phase_controller_inst1_state_4;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.time_passed11 ;
    wire \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.hc_time_passed ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.N_279 ;
    wire \phase_controller_inst1.stoper_tr.N_262 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_335_i_g ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_reg3lto19_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_18_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_18_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_18_17_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_18_18_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_337_i ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_18_19_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_18_20_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire bfn_18_21_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_reg3lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_320_4 ;
    wire \delay_measurement_inst.delay_tr_timer.N_320_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.N_328 ;
    wire \delay_measurement_inst.delay_tr_timer.N_331_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ;
    wire \delay_measurement_inst.delay_tr_timer.N_321_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.N_331 ;
    wire \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14 ;
    wire \delay_measurement_inst.delay_tr_reg3lto14 ;
    wire measured_delay_tr_14;
    wire \delay_measurement_inst.delay_tr_reg3lto15 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ;
    wire measured_delay_tr_15;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire measured_delay_tr_1;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire measured_delay_tr_5;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire measured_delay_tr_3;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire measured_delay_tr_8;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire measured_delay_tr_7;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire measured_delay_tr_13;
    wire \delay_measurement_inst.delay_tr_reg3lto6 ;
    wire measured_delay_tr_6;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire measured_delay_tr_4;
    wire \delay_measurement_inst.N_324 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire measured_delay_tr_2;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.N_301 ;
    wire measured_delay_tr_11;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire measured_delay_tr_18;
    wire measured_delay_tr_17;
    wire measured_delay_tr_16;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_i ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.N_358 ;
    wire measured_delay_tr_19;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__20819),
            .RESETB(N__35880),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__23099),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__23089),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__20529,N__20557,N__20530,N__20558,N__20531,N__18716,N__18740,N__18779,N__18692,N__18758,N__19525,N__19551,N__18643,N__18631,N__18655}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__23095,N__23092,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__23090,N__23094,N__23091,N__23093}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__23064),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__23057),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64}),
            .ADDSUBBOT(),
            .A({dangling_wire_65,N__20612,N__20605,N__20610,N__20604,N__20611,N__20603,N__20613,N__20600,N__20606,N__20599,N__20607,N__20601,N__20608,N__20602,N__20609}),
            .C({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .B({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__23063,N__23060,dangling_wire_89,dangling_wire_90,dangling_wire_91,N__23058,N__23062,N__23059,N__23061}),
            .OHOLDTOP(),
            .O({dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__48678),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__48680),
            .DIN(N__48679),
            .DOUT(N__48678),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__48680),
            .PADOUT(N__48679),
            .PADIN(N__48678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__48669),
            .DIN(N__48668),
            .DOUT(N__48667),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__48669),
            .PADOUT(N__48668),
            .PADIN(N__48667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__48660),
            .DIN(N__48659),
            .DOUT(N__48658),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__48660),
            .PADOUT(N__48659),
            .PADIN(N__48658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__48651),
            .DIN(N__48650),
            .DOUT(N__48649),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__48651),
            .PADOUT(N__48650),
            .PADIN(N__48649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__48642),
            .DIN(N__48641),
            .DOUT(N__48640),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__48642),
            .PADOUT(N__48641),
            .PADIN(N__48640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__48633),
            .DIN(N__48632),
            .DOUT(N__48631),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__48633),
            .PADOUT(N__48632),
            .PADIN(N__48631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34073),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__48624),
            .DIN(N__48623),
            .DOUT(N__48622),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__48624),
            .PADOUT(N__48623),
            .PADIN(N__48622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__48615),
            .DIN(N__48614),
            .DOUT(N__48613),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__48615),
            .PADOUT(N__48614),
            .PADIN(N__48613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__48606),
            .DIN(N__48605),
            .DOUT(N__48604),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__48606),
            .PADOUT(N__48605),
            .PADIN(N__48604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__48597),
            .DIN(N__48596),
            .DOUT(N__48595),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__48597),
            .PADOUT(N__48596),
            .PADIN(N__48595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32327),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__48588),
            .DIN(N__48587),
            .DOUT(N__48586),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__48588),
            .PADOUT(N__48587),
            .PADIN(N__48586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33641),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__48579),
            .DIN(N__48578),
            .DOUT(N__48577),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__48579),
            .PADOUT(N__48578),
            .PADIN(N__48577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__48570),
            .DIN(N__48569),
            .DOUT(N__48568),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__48570),
            .PADOUT(N__48569),
            .PADIN(N__48568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11621 (
            .O(N__48551),
            .I(N__48547));
    InMux I__11620 (
            .O(N__48550),
            .I(N__48544));
    LocalMux I__11619 (
            .O(N__48547),
            .I(N__48538));
    LocalMux I__11618 (
            .O(N__48544),
            .I(N__48538));
    InMux I__11617 (
            .O(N__48543),
            .I(N__48535));
    Span4Mux_v I__11616 (
            .O(N__48538),
            .I(N__48532));
    LocalMux I__11615 (
            .O(N__48535),
            .I(N__48529));
    Odrv4 I__11614 (
            .O(N__48532),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    Odrv4 I__11613 (
            .O(N__48529),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__11612 (
            .O(N__48524),
            .I(N__48521));
    LocalMux I__11611 (
            .O(N__48521),
            .I(N__48517));
    InMux I__11610 (
            .O(N__48520),
            .I(N__48514));
    Span4Mux_v I__11609 (
            .O(N__48517),
            .I(N__48509));
    LocalMux I__11608 (
            .O(N__48514),
            .I(N__48509));
    Odrv4 I__11607 (
            .O(N__48509),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__11606 (
            .O(N__48506),
            .I(N__48499));
    InMux I__11605 (
            .O(N__48505),
            .I(N__48499));
    InMux I__11604 (
            .O(N__48504),
            .I(N__48496));
    LocalMux I__11603 (
            .O(N__48499),
            .I(N__48491));
    LocalMux I__11602 (
            .O(N__48496),
            .I(N__48488));
    InMux I__11601 (
            .O(N__48495),
            .I(N__48485));
    InMux I__11600 (
            .O(N__48494),
            .I(N__48482));
    Span4Mux_h I__11599 (
            .O(N__48491),
            .I(N__48479));
    Span4Mux_h I__11598 (
            .O(N__48488),
            .I(N__48472));
    LocalMux I__11597 (
            .O(N__48485),
            .I(N__48472));
    LocalMux I__11596 (
            .O(N__48482),
            .I(N__48472));
    Odrv4 I__11595 (
            .O(N__48479),
            .I(\delay_measurement_inst.N_301 ));
    Odrv4 I__11594 (
            .O(N__48472),
            .I(\delay_measurement_inst.N_301 ));
    InMux I__11593 (
            .O(N__48467),
            .I(N__48463));
    InMux I__11592 (
            .O(N__48466),
            .I(N__48460));
    LocalMux I__11591 (
            .O(N__48463),
            .I(N__48454));
    LocalMux I__11590 (
            .O(N__48460),
            .I(N__48454));
    InMux I__11589 (
            .O(N__48459),
            .I(N__48451));
    Span12Mux_s10_v I__11588 (
            .O(N__48454),
            .I(N__48446));
    LocalMux I__11587 (
            .O(N__48451),
            .I(N__48446));
    Odrv12 I__11586 (
            .O(N__48446),
            .I(measured_delay_tr_11));
    InMux I__11585 (
            .O(N__48443),
            .I(N__48439));
    InMux I__11584 (
            .O(N__48442),
            .I(N__48435));
    LocalMux I__11583 (
            .O(N__48439),
            .I(N__48432));
    InMux I__11582 (
            .O(N__48438),
            .I(N__48429));
    LocalMux I__11581 (
            .O(N__48435),
            .I(N__48426));
    Span4Mux_v I__11580 (
            .O(N__48432),
            .I(N__48423));
    LocalMux I__11579 (
            .O(N__48429),
            .I(N__48420));
    Span4Mux_h I__11578 (
            .O(N__48426),
            .I(N__48417));
    Odrv4 I__11577 (
            .O(N__48423),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv12 I__11576 (
            .O(N__48420),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__11575 (
            .O(N__48417),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__11574 (
            .O(N__48410),
            .I(N__48406));
    InMux I__11573 (
            .O(N__48409),
            .I(N__48403));
    LocalMux I__11572 (
            .O(N__48406),
            .I(N__48397));
    LocalMux I__11571 (
            .O(N__48403),
            .I(N__48397));
    InMux I__11570 (
            .O(N__48402),
            .I(N__48394));
    Span4Mux_v I__11569 (
            .O(N__48397),
            .I(N__48389));
    LocalMux I__11568 (
            .O(N__48394),
            .I(N__48389));
    Span4Mux_h I__11567 (
            .O(N__48389),
            .I(N__48385));
    InMux I__11566 (
            .O(N__48388),
            .I(N__48382));
    Odrv4 I__11565 (
            .O(N__48385),
            .I(measured_delay_tr_18));
    LocalMux I__11564 (
            .O(N__48382),
            .I(measured_delay_tr_18));
    InMux I__11563 (
            .O(N__48377),
            .I(N__48374));
    LocalMux I__11562 (
            .O(N__48374),
            .I(N__48370));
    InMux I__11561 (
            .O(N__48373),
            .I(N__48367));
    Span4Mux_v I__11560 (
            .O(N__48370),
            .I(N__48361));
    LocalMux I__11559 (
            .O(N__48367),
            .I(N__48361));
    InMux I__11558 (
            .O(N__48366),
            .I(N__48358));
    Span4Mux_h I__11557 (
            .O(N__48361),
            .I(N__48352));
    LocalMux I__11556 (
            .O(N__48358),
            .I(N__48352));
    InMux I__11555 (
            .O(N__48357),
            .I(N__48349));
    Span4Mux_v I__11554 (
            .O(N__48352),
            .I(N__48346));
    LocalMux I__11553 (
            .O(N__48349),
            .I(N__48343));
    Odrv4 I__11552 (
            .O(N__48346),
            .I(measured_delay_tr_17));
    Odrv4 I__11551 (
            .O(N__48343),
            .I(measured_delay_tr_17));
    InMux I__11550 (
            .O(N__48338),
            .I(N__48335));
    LocalMux I__11549 (
            .O(N__48335),
            .I(N__48331));
    InMux I__11548 (
            .O(N__48334),
            .I(N__48328));
    Span4Mux_v I__11547 (
            .O(N__48331),
            .I(N__48322));
    LocalMux I__11546 (
            .O(N__48328),
            .I(N__48322));
    InMux I__11545 (
            .O(N__48327),
            .I(N__48319));
    Span4Mux_h I__11544 (
            .O(N__48322),
            .I(N__48313));
    LocalMux I__11543 (
            .O(N__48319),
            .I(N__48313));
    InMux I__11542 (
            .O(N__48318),
            .I(N__48310));
    Span4Mux_h I__11541 (
            .O(N__48313),
            .I(N__48307));
    LocalMux I__11540 (
            .O(N__48310),
            .I(N__48304));
    Odrv4 I__11539 (
            .O(N__48307),
            .I(measured_delay_tr_16));
    Odrv4 I__11538 (
            .O(N__48304),
            .I(measured_delay_tr_16));
    InMux I__11537 (
            .O(N__48299),
            .I(N__48296));
    LocalMux I__11536 (
            .O(N__48296),
            .I(N__48293));
    Odrv4 I__11535 (
            .O(N__48293),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ));
    InMux I__11534 (
            .O(N__48290),
            .I(N__48287));
    LocalMux I__11533 (
            .O(N__48287),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_i ));
    CascadeMux I__11532 (
            .O(N__48284),
            .I(N__48275));
    CascadeMux I__11531 (
            .O(N__48283),
            .I(N__48270));
    CascadeMux I__11530 (
            .O(N__48282),
            .I(N__48267));
    CascadeMux I__11529 (
            .O(N__48281),
            .I(N__48262));
    InMux I__11528 (
            .O(N__48280),
            .I(N__48254));
    InMux I__11527 (
            .O(N__48279),
            .I(N__48247));
    InMux I__11526 (
            .O(N__48278),
            .I(N__48247));
    InMux I__11525 (
            .O(N__48275),
            .I(N__48240));
    InMux I__11524 (
            .O(N__48274),
            .I(N__48240));
    InMux I__11523 (
            .O(N__48273),
            .I(N__48240));
    InMux I__11522 (
            .O(N__48270),
            .I(N__48231));
    InMux I__11521 (
            .O(N__48267),
            .I(N__48231));
    InMux I__11520 (
            .O(N__48266),
            .I(N__48231));
    InMux I__11519 (
            .O(N__48265),
            .I(N__48231));
    InMux I__11518 (
            .O(N__48262),
            .I(N__48228));
    InMux I__11517 (
            .O(N__48261),
            .I(N__48223));
    InMux I__11516 (
            .O(N__48260),
            .I(N__48223));
    CascadeMux I__11515 (
            .O(N__48259),
            .I(N__48220));
    CascadeMux I__11514 (
            .O(N__48258),
            .I(N__48217));
    CascadeMux I__11513 (
            .O(N__48257),
            .I(N__48212));
    LocalMux I__11512 (
            .O(N__48254),
            .I(N__48208));
    InMux I__11511 (
            .O(N__48253),
            .I(N__48203));
    InMux I__11510 (
            .O(N__48252),
            .I(N__48203));
    LocalMux I__11509 (
            .O(N__48247),
            .I(N__48196));
    LocalMux I__11508 (
            .O(N__48240),
            .I(N__48196));
    LocalMux I__11507 (
            .O(N__48231),
            .I(N__48196));
    LocalMux I__11506 (
            .O(N__48228),
            .I(N__48191));
    LocalMux I__11505 (
            .O(N__48223),
            .I(N__48191));
    InMux I__11504 (
            .O(N__48220),
            .I(N__48178));
    InMux I__11503 (
            .O(N__48217),
            .I(N__48178));
    InMux I__11502 (
            .O(N__48216),
            .I(N__48178));
    InMux I__11501 (
            .O(N__48215),
            .I(N__48178));
    InMux I__11500 (
            .O(N__48212),
            .I(N__48178));
    InMux I__11499 (
            .O(N__48211),
            .I(N__48178));
    Span4Mux_v I__11498 (
            .O(N__48208),
            .I(N__48173));
    LocalMux I__11497 (
            .O(N__48203),
            .I(N__48173));
    Span4Mux_v I__11496 (
            .O(N__48196),
            .I(N__48168));
    Span4Mux_v I__11495 (
            .O(N__48191),
            .I(N__48168));
    LocalMux I__11494 (
            .O(N__48178),
            .I(N__48165));
    Span4Mux_h I__11493 (
            .O(N__48173),
            .I(N__48162));
    Odrv4 I__11492 (
            .O(N__48168),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv12 I__11491 (
            .O(N__48165),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__11490 (
            .O(N__48162),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    InMux I__11489 (
            .O(N__48155),
            .I(N__48151));
    InMux I__11488 (
            .O(N__48154),
            .I(N__48148));
    LocalMux I__11487 (
            .O(N__48151),
            .I(N__48144));
    LocalMux I__11486 (
            .O(N__48148),
            .I(N__48141));
    CascadeMux I__11485 (
            .O(N__48147),
            .I(N__48138));
    Span4Mux_v I__11484 (
            .O(N__48144),
            .I(N__48133));
    Span4Mux_v I__11483 (
            .O(N__48141),
            .I(N__48133));
    InMux I__11482 (
            .O(N__48138),
            .I(N__48130));
    Sp12to4 I__11481 (
            .O(N__48133),
            .I(N__48125));
    LocalMux I__11480 (
            .O(N__48130),
            .I(N__48125));
    Odrv12 I__11479 (
            .O(N__48125),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__11478 (
            .O(N__48122),
            .I(N__48114));
    InMux I__11477 (
            .O(N__48121),
            .I(N__48114));
    InMux I__11476 (
            .O(N__48120),
            .I(N__48111));
    InMux I__11475 (
            .O(N__48119),
            .I(N__48108));
    LocalMux I__11474 (
            .O(N__48114),
            .I(N__48103));
    LocalMux I__11473 (
            .O(N__48111),
            .I(N__48100));
    LocalMux I__11472 (
            .O(N__48108),
            .I(N__48097));
    InMux I__11471 (
            .O(N__48107),
            .I(N__48092));
    InMux I__11470 (
            .O(N__48106),
            .I(N__48092));
    Span4Mux_v I__11469 (
            .O(N__48103),
            .I(N__48081));
    Span4Mux_h I__11468 (
            .O(N__48100),
            .I(N__48081));
    Span4Mux_v I__11467 (
            .O(N__48097),
            .I(N__48081));
    LocalMux I__11466 (
            .O(N__48092),
            .I(N__48081));
    InMux I__11465 (
            .O(N__48091),
            .I(N__48075));
    InMux I__11464 (
            .O(N__48090),
            .I(N__48075));
    Span4Mux_h I__11463 (
            .O(N__48081),
            .I(N__48072));
    InMux I__11462 (
            .O(N__48080),
            .I(N__48069));
    LocalMux I__11461 (
            .O(N__48075),
            .I(N__48066));
    Odrv4 I__11460 (
            .O(N__48072),
            .I(\delay_measurement_inst.N_358 ));
    LocalMux I__11459 (
            .O(N__48069),
            .I(\delay_measurement_inst.N_358 ));
    Odrv12 I__11458 (
            .O(N__48066),
            .I(\delay_measurement_inst.N_358 ));
    InMux I__11457 (
            .O(N__48059),
            .I(N__48056));
    LocalMux I__11456 (
            .O(N__48056),
            .I(N__48051));
    CascadeMux I__11455 (
            .O(N__48055),
            .I(N__48048));
    InMux I__11454 (
            .O(N__48054),
            .I(N__48045));
    Span4Mux_v I__11453 (
            .O(N__48051),
            .I(N__48041));
    InMux I__11452 (
            .O(N__48048),
            .I(N__48038));
    LocalMux I__11451 (
            .O(N__48045),
            .I(N__48035));
    CascadeMux I__11450 (
            .O(N__48044),
            .I(N__48032));
    Span4Mux_h I__11449 (
            .O(N__48041),
            .I(N__48027));
    LocalMux I__11448 (
            .O(N__48038),
            .I(N__48027));
    Span4Mux_v I__11447 (
            .O(N__48035),
            .I(N__48024));
    InMux I__11446 (
            .O(N__48032),
            .I(N__48021));
    Span4Mux_v I__11445 (
            .O(N__48027),
            .I(N__48018));
    Span4Mux_h I__11444 (
            .O(N__48024),
            .I(N__48013));
    LocalMux I__11443 (
            .O(N__48021),
            .I(N__48013));
    Odrv4 I__11442 (
            .O(N__48018),
            .I(measured_delay_tr_19));
    Odrv4 I__11441 (
            .O(N__48013),
            .I(measured_delay_tr_19));
    ClkMux I__11440 (
            .O(N__48008),
            .I(N__47522));
    ClkMux I__11439 (
            .O(N__48007),
            .I(N__47522));
    ClkMux I__11438 (
            .O(N__48006),
            .I(N__47522));
    ClkMux I__11437 (
            .O(N__48005),
            .I(N__47522));
    ClkMux I__11436 (
            .O(N__48004),
            .I(N__47522));
    ClkMux I__11435 (
            .O(N__48003),
            .I(N__47522));
    ClkMux I__11434 (
            .O(N__48002),
            .I(N__47522));
    ClkMux I__11433 (
            .O(N__48001),
            .I(N__47522));
    ClkMux I__11432 (
            .O(N__48000),
            .I(N__47522));
    ClkMux I__11431 (
            .O(N__47999),
            .I(N__47522));
    ClkMux I__11430 (
            .O(N__47998),
            .I(N__47522));
    ClkMux I__11429 (
            .O(N__47997),
            .I(N__47522));
    ClkMux I__11428 (
            .O(N__47996),
            .I(N__47522));
    ClkMux I__11427 (
            .O(N__47995),
            .I(N__47522));
    ClkMux I__11426 (
            .O(N__47994),
            .I(N__47522));
    ClkMux I__11425 (
            .O(N__47993),
            .I(N__47522));
    ClkMux I__11424 (
            .O(N__47992),
            .I(N__47522));
    ClkMux I__11423 (
            .O(N__47991),
            .I(N__47522));
    ClkMux I__11422 (
            .O(N__47990),
            .I(N__47522));
    ClkMux I__11421 (
            .O(N__47989),
            .I(N__47522));
    ClkMux I__11420 (
            .O(N__47988),
            .I(N__47522));
    ClkMux I__11419 (
            .O(N__47987),
            .I(N__47522));
    ClkMux I__11418 (
            .O(N__47986),
            .I(N__47522));
    ClkMux I__11417 (
            .O(N__47985),
            .I(N__47522));
    ClkMux I__11416 (
            .O(N__47984),
            .I(N__47522));
    ClkMux I__11415 (
            .O(N__47983),
            .I(N__47522));
    ClkMux I__11414 (
            .O(N__47982),
            .I(N__47522));
    ClkMux I__11413 (
            .O(N__47981),
            .I(N__47522));
    ClkMux I__11412 (
            .O(N__47980),
            .I(N__47522));
    ClkMux I__11411 (
            .O(N__47979),
            .I(N__47522));
    ClkMux I__11410 (
            .O(N__47978),
            .I(N__47522));
    ClkMux I__11409 (
            .O(N__47977),
            .I(N__47522));
    ClkMux I__11408 (
            .O(N__47976),
            .I(N__47522));
    ClkMux I__11407 (
            .O(N__47975),
            .I(N__47522));
    ClkMux I__11406 (
            .O(N__47974),
            .I(N__47522));
    ClkMux I__11405 (
            .O(N__47973),
            .I(N__47522));
    ClkMux I__11404 (
            .O(N__47972),
            .I(N__47522));
    ClkMux I__11403 (
            .O(N__47971),
            .I(N__47522));
    ClkMux I__11402 (
            .O(N__47970),
            .I(N__47522));
    ClkMux I__11401 (
            .O(N__47969),
            .I(N__47522));
    ClkMux I__11400 (
            .O(N__47968),
            .I(N__47522));
    ClkMux I__11399 (
            .O(N__47967),
            .I(N__47522));
    ClkMux I__11398 (
            .O(N__47966),
            .I(N__47522));
    ClkMux I__11397 (
            .O(N__47965),
            .I(N__47522));
    ClkMux I__11396 (
            .O(N__47964),
            .I(N__47522));
    ClkMux I__11395 (
            .O(N__47963),
            .I(N__47522));
    ClkMux I__11394 (
            .O(N__47962),
            .I(N__47522));
    ClkMux I__11393 (
            .O(N__47961),
            .I(N__47522));
    ClkMux I__11392 (
            .O(N__47960),
            .I(N__47522));
    ClkMux I__11391 (
            .O(N__47959),
            .I(N__47522));
    ClkMux I__11390 (
            .O(N__47958),
            .I(N__47522));
    ClkMux I__11389 (
            .O(N__47957),
            .I(N__47522));
    ClkMux I__11388 (
            .O(N__47956),
            .I(N__47522));
    ClkMux I__11387 (
            .O(N__47955),
            .I(N__47522));
    ClkMux I__11386 (
            .O(N__47954),
            .I(N__47522));
    ClkMux I__11385 (
            .O(N__47953),
            .I(N__47522));
    ClkMux I__11384 (
            .O(N__47952),
            .I(N__47522));
    ClkMux I__11383 (
            .O(N__47951),
            .I(N__47522));
    ClkMux I__11382 (
            .O(N__47950),
            .I(N__47522));
    ClkMux I__11381 (
            .O(N__47949),
            .I(N__47522));
    ClkMux I__11380 (
            .O(N__47948),
            .I(N__47522));
    ClkMux I__11379 (
            .O(N__47947),
            .I(N__47522));
    ClkMux I__11378 (
            .O(N__47946),
            .I(N__47522));
    ClkMux I__11377 (
            .O(N__47945),
            .I(N__47522));
    ClkMux I__11376 (
            .O(N__47944),
            .I(N__47522));
    ClkMux I__11375 (
            .O(N__47943),
            .I(N__47522));
    ClkMux I__11374 (
            .O(N__47942),
            .I(N__47522));
    ClkMux I__11373 (
            .O(N__47941),
            .I(N__47522));
    ClkMux I__11372 (
            .O(N__47940),
            .I(N__47522));
    ClkMux I__11371 (
            .O(N__47939),
            .I(N__47522));
    ClkMux I__11370 (
            .O(N__47938),
            .I(N__47522));
    ClkMux I__11369 (
            .O(N__47937),
            .I(N__47522));
    ClkMux I__11368 (
            .O(N__47936),
            .I(N__47522));
    ClkMux I__11367 (
            .O(N__47935),
            .I(N__47522));
    ClkMux I__11366 (
            .O(N__47934),
            .I(N__47522));
    ClkMux I__11365 (
            .O(N__47933),
            .I(N__47522));
    ClkMux I__11364 (
            .O(N__47932),
            .I(N__47522));
    ClkMux I__11363 (
            .O(N__47931),
            .I(N__47522));
    ClkMux I__11362 (
            .O(N__47930),
            .I(N__47522));
    ClkMux I__11361 (
            .O(N__47929),
            .I(N__47522));
    ClkMux I__11360 (
            .O(N__47928),
            .I(N__47522));
    ClkMux I__11359 (
            .O(N__47927),
            .I(N__47522));
    ClkMux I__11358 (
            .O(N__47926),
            .I(N__47522));
    ClkMux I__11357 (
            .O(N__47925),
            .I(N__47522));
    ClkMux I__11356 (
            .O(N__47924),
            .I(N__47522));
    ClkMux I__11355 (
            .O(N__47923),
            .I(N__47522));
    ClkMux I__11354 (
            .O(N__47922),
            .I(N__47522));
    ClkMux I__11353 (
            .O(N__47921),
            .I(N__47522));
    ClkMux I__11352 (
            .O(N__47920),
            .I(N__47522));
    ClkMux I__11351 (
            .O(N__47919),
            .I(N__47522));
    ClkMux I__11350 (
            .O(N__47918),
            .I(N__47522));
    ClkMux I__11349 (
            .O(N__47917),
            .I(N__47522));
    ClkMux I__11348 (
            .O(N__47916),
            .I(N__47522));
    ClkMux I__11347 (
            .O(N__47915),
            .I(N__47522));
    ClkMux I__11346 (
            .O(N__47914),
            .I(N__47522));
    ClkMux I__11345 (
            .O(N__47913),
            .I(N__47522));
    ClkMux I__11344 (
            .O(N__47912),
            .I(N__47522));
    ClkMux I__11343 (
            .O(N__47911),
            .I(N__47522));
    ClkMux I__11342 (
            .O(N__47910),
            .I(N__47522));
    ClkMux I__11341 (
            .O(N__47909),
            .I(N__47522));
    ClkMux I__11340 (
            .O(N__47908),
            .I(N__47522));
    ClkMux I__11339 (
            .O(N__47907),
            .I(N__47522));
    ClkMux I__11338 (
            .O(N__47906),
            .I(N__47522));
    ClkMux I__11337 (
            .O(N__47905),
            .I(N__47522));
    ClkMux I__11336 (
            .O(N__47904),
            .I(N__47522));
    ClkMux I__11335 (
            .O(N__47903),
            .I(N__47522));
    ClkMux I__11334 (
            .O(N__47902),
            .I(N__47522));
    ClkMux I__11333 (
            .O(N__47901),
            .I(N__47522));
    ClkMux I__11332 (
            .O(N__47900),
            .I(N__47522));
    ClkMux I__11331 (
            .O(N__47899),
            .I(N__47522));
    ClkMux I__11330 (
            .O(N__47898),
            .I(N__47522));
    ClkMux I__11329 (
            .O(N__47897),
            .I(N__47522));
    ClkMux I__11328 (
            .O(N__47896),
            .I(N__47522));
    ClkMux I__11327 (
            .O(N__47895),
            .I(N__47522));
    ClkMux I__11326 (
            .O(N__47894),
            .I(N__47522));
    ClkMux I__11325 (
            .O(N__47893),
            .I(N__47522));
    ClkMux I__11324 (
            .O(N__47892),
            .I(N__47522));
    ClkMux I__11323 (
            .O(N__47891),
            .I(N__47522));
    ClkMux I__11322 (
            .O(N__47890),
            .I(N__47522));
    ClkMux I__11321 (
            .O(N__47889),
            .I(N__47522));
    ClkMux I__11320 (
            .O(N__47888),
            .I(N__47522));
    ClkMux I__11319 (
            .O(N__47887),
            .I(N__47522));
    ClkMux I__11318 (
            .O(N__47886),
            .I(N__47522));
    ClkMux I__11317 (
            .O(N__47885),
            .I(N__47522));
    ClkMux I__11316 (
            .O(N__47884),
            .I(N__47522));
    ClkMux I__11315 (
            .O(N__47883),
            .I(N__47522));
    ClkMux I__11314 (
            .O(N__47882),
            .I(N__47522));
    ClkMux I__11313 (
            .O(N__47881),
            .I(N__47522));
    ClkMux I__11312 (
            .O(N__47880),
            .I(N__47522));
    ClkMux I__11311 (
            .O(N__47879),
            .I(N__47522));
    ClkMux I__11310 (
            .O(N__47878),
            .I(N__47522));
    ClkMux I__11309 (
            .O(N__47877),
            .I(N__47522));
    ClkMux I__11308 (
            .O(N__47876),
            .I(N__47522));
    ClkMux I__11307 (
            .O(N__47875),
            .I(N__47522));
    ClkMux I__11306 (
            .O(N__47874),
            .I(N__47522));
    ClkMux I__11305 (
            .O(N__47873),
            .I(N__47522));
    ClkMux I__11304 (
            .O(N__47872),
            .I(N__47522));
    ClkMux I__11303 (
            .O(N__47871),
            .I(N__47522));
    ClkMux I__11302 (
            .O(N__47870),
            .I(N__47522));
    ClkMux I__11301 (
            .O(N__47869),
            .I(N__47522));
    ClkMux I__11300 (
            .O(N__47868),
            .I(N__47522));
    ClkMux I__11299 (
            .O(N__47867),
            .I(N__47522));
    ClkMux I__11298 (
            .O(N__47866),
            .I(N__47522));
    ClkMux I__11297 (
            .O(N__47865),
            .I(N__47522));
    ClkMux I__11296 (
            .O(N__47864),
            .I(N__47522));
    ClkMux I__11295 (
            .O(N__47863),
            .I(N__47522));
    ClkMux I__11294 (
            .O(N__47862),
            .I(N__47522));
    ClkMux I__11293 (
            .O(N__47861),
            .I(N__47522));
    ClkMux I__11292 (
            .O(N__47860),
            .I(N__47522));
    ClkMux I__11291 (
            .O(N__47859),
            .I(N__47522));
    ClkMux I__11290 (
            .O(N__47858),
            .I(N__47522));
    ClkMux I__11289 (
            .O(N__47857),
            .I(N__47522));
    ClkMux I__11288 (
            .O(N__47856),
            .I(N__47522));
    ClkMux I__11287 (
            .O(N__47855),
            .I(N__47522));
    ClkMux I__11286 (
            .O(N__47854),
            .I(N__47522));
    ClkMux I__11285 (
            .O(N__47853),
            .I(N__47522));
    ClkMux I__11284 (
            .O(N__47852),
            .I(N__47522));
    ClkMux I__11283 (
            .O(N__47851),
            .I(N__47522));
    ClkMux I__11282 (
            .O(N__47850),
            .I(N__47522));
    ClkMux I__11281 (
            .O(N__47849),
            .I(N__47522));
    ClkMux I__11280 (
            .O(N__47848),
            .I(N__47522));
    ClkMux I__11279 (
            .O(N__47847),
            .I(N__47522));
    GlobalMux I__11278 (
            .O(N__47522),
            .I(clk_100mhz_0));
    CEMux I__11277 (
            .O(N__47519),
            .I(N__47515));
    CEMux I__11276 (
            .O(N__47518),
            .I(N__47512));
    LocalMux I__11275 (
            .O(N__47515),
            .I(N__47508));
    LocalMux I__11274 (
            .O(N__47512),
            .I(N__47505));
    CEMux I__11273 (
            .O(N__47511),
            .I(N__47502));
    Span4Mux_v I__11272 (
            .O(N__47508),
            .I(N__47499));
    Span4Mux_v I__11271 (
            .O(N__47505),
            .I(N__47496));
    LocalMux I__11270 (
            .O(N__47502),
            .I(N__47493));
    Span4Mux_h I__11269 (
            .O(N__47499),
            .I(N__47483));
    Span4Mux_h I__11268 (
            .O(N__47496),
            .I(N__47483));
    Span4Mux_v I__11267 (
            .O(N__47493),
            .I(N__47483));
    CEMux I__11266 (
            .O(N__47492),
            .I(N__47480));
    CEMux I__11265 (
            .O(N__47491),
            .I(N__47477));
    CEMux I__11264 (
            .O(N__47490),
            .I(N__47474));
    Odrv4 I__11263 (
            .O(N__47483),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__11262 (
            .O(N__47480),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__11261 (
            .O(N__47477),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__11260 (
            .O(N__47474),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    CascadeMux I__11259 (
            .O(N__47465),
            .I(N__47456));
    CascadeMux I__11258 (
            .O(N__47464),
            .I(N__47453));
    InMux I__11257 (
            .O(N__47463),
            .I(N__47450));
    InMux I__11256 (
            .O(N__47462),
            .I(N__47447));
    InMux I__11255 (
            .O(N__47461),
            .I(N__47444));
    InMux I__11254 (
            .O(N__47460),
            .I(N__47441));
    InMux I__11253 (
            .O(N__47459),
            .I(N__47438));
    InMux I__11252 (
            .O(N__47456),
            .I(N__47435));
    InMux I__11251 (
            .O(N__47453),
            .I(N__47432));
    LocalMux I__11250 (
            .O(N__47450),
            .I(N__47429));
    LocalMux I__11249 (
            .O(N__47447),
            .I(N__47426));
    LocalMux I__11248 (
            .O(N__47444),
            .I(N__47423));
    LocalMux I__11247 (
            .O(N__47441),
            .I(N__47418));
    LocalMux I__11246 (
            .O(N__47438),
            .I(N__47332));
    LocalMux I__11245 (
            .O(N__47435),
            .I(N__47283));
    LocalMux I__11244 (
            .O(N__47432),
            .I(N__47280));
    Glb2LocalMux I__11243 (
            .O(N__47429),
            .I(N__46979));
    Glb2LocalMux I__11242 (
            .O(N__47426),
            .I(N__46979));
    Glb2LocalMux I__11241 (
            .O(N__47423),
            .I(N__46979));
    SRMux I__11240 (
            .O(N__47422),
            .I(N__46979));
    SRMux I__11239 (
            .O(N__47421),
            .I(N__46979));
    Glb2LocalMux I__11238 (
            .O(N__47418),
            .I(N__46979));
    SRMux I__11237 (
            .O(N__47417),
            .I(N__46979));
    SRMux I__11236 (
            .O(N__47416),
            .I(N__46979));
    SRMux I__11235 (
            .O(N__47415),
            .I(N__46979));
    SRMux I__11234 (
            .O(N__47414),
            .I(N__46979));
    SRMux I__11233 (
            .O(N__47413),
            .I(N__46979));
    SRMux I__11232 (
            .O(N__47412),
            .I(N__46979));
    SRMux I__11231 (
            .O(N__47411),
            .I(N__46979));
    SRMux I__11230 (
            .O(N__47410),
            .I(N__46979));
    SRMux I__11229 (
            .O(N__47409),
            .I(N__46979));
    SRMux I__11228 (
            .O(N__47408),
            .I(N__46979));
    SRMux I__11227 (
            .O(N__47407),
            .I(N__46979));
    SRMux I__11226 (
            .O(N__47406),
            .I(N__46979));
    SRMux I__11225 (
            .O(N__47405),
            .I(N__46979));
    SRMux I__11224 (
            .O(N__47404),
            .I(N__46979));
    SRMux I__11223 (
            .O(N__47403),
            .I(N__46979));
    SRMux I__11222 (
            .O(N__47402),
            .I(N__46979));
    SRMux I__11221 (
            .O(N__47401),
            .I(N__46979));
    SRMux I__11220 (
            .O(N__47400),
            .I(N__46979));
    SRMux I__11219 (
            .O(N__47399),
            .I(N__46979));
    SRMux I__11218 (
            .O(N__47398),
            .I(N__46979));
    SRMux I__11217 (
            .O(N__47397),
            .I(N__46979));
    SRMux I__11216 (
            .O(N__47396),
            .I(N__46979));
    SRMux I__11215 (
            .O(N__47395),
            .I(N__46979));
    SRMux I__11214 (
            .O(N__47394),
            .I(N__46979));
    SRMux I__11213 (
            .O(N__47393),
            .I(N__46979));
    SRMux I__11212 (
            .O(N__47392),
            .I(N__46979));
    SRMux I__11211 (
            .O(N__47391),
            .I(N__46979));
    SRMux I__11210 (
            .O(N__47390),
            .I(N__46979));
    SRMux I__11209 (
            .O(N__47389),
            .I(N__46979));
    SRMux I__11208 (
            .O(N__47388),
            .I(N__46979));
    SRMux I__11207 (
            .O(N__47387),
            .I(N__46979));
    SRMux I__11206 (
            .O(N__47386),
            .I(N__46979));
    SRMux I__11205 (
            .O(N__47385),
            .I(N__46979));
    SRMux I__11204 (
            .O(N__47384),
            .I(N__46979));
    SRMux I__11203 (
            .O(N__47383),
            .I(N__46979));
    SRMux I__11202 (
            .O(N__47382),
            .I(N__46979));
    SRMux I__11201 (
            .O(N__47381),
            .I(N__46979));
    SRMux I__11200 (
            .O(N__47380),
            .I(N__46979));
    SRMux I__11199 (
            .O(N__47379),
            .I(N__46979));
    SRMux I__11198 (
            .O(N__47378),
            .I(N__46979));
    SRMux I__11197 (
            .O(N__47377),
            .I(N__46979));
    SRMux I__11196 (
            .O(N__47376),
            .I(N__46979));
    SRMux I__11195 (
            .O(N__47375),
            .I(N__46979));
    SRMux I__11194 (
            .O(N__47374),
            .I(N__46979));
    SRMux I__11193 (
            .O(N__47373),
            .I(N__46979));
    SRMux I__11192 (
            .O(N__47372),
            .I(N__46979));
    SRMux I__11191 (
            .O(N__47371),
            .I(N__46979));
    SRMux I__11190 (
            .O(N__47370),
            .I(N__46979));
    SRMux I__11189 (
            .O(N__47369),
            .I(N__46979));
    SRMux I__11188 (
            .O(N__47368),
            .I(N__46979));
    SRMux I__11187 (
            .O(N__47367),
            .I(N__46979));
    SRMux I__11186 (
            .O(N__47366),
            .I(N__46979));
    SRMux I__11185 (
            .O(N__47365),
            .I(N__46979));
    SRMux I__11184 (
            .O(N__47364),
            .I(N__46979));
    SRMux I__11183 (
            .O(N__47363),
            .I(N__46979));
    SRMux I__11182 (
            .O(N__47362),
            .I(N__46979));
    SRMux I__11181 (
            .O(N__47361),
            .I(N__46979));
    SRMux I__11180 (
            .O(N__47360),
            .I(N__46979));
    SRMux I__11179 (
            .O(N__47359),
            .I(N__46979));
    SRMux I__11178 (
            .O(N__47358),
            .I(N__46979));
    SRMux I__11177 (
            .O(N__47357),
            .I(N__46979));
    SRMux I__11176 (
            .O(N__47356),
            .I(N__46979));
    SRMux I__11175 (
            .O(N__47355),
            .I(N__46979));
    SRMux I__11174 (
            .O(N__47354),
            .I(N__46979));
    SRMux I__11173 (
            .O(N__47353),
            .I(N__46979));
    SRMux I__11172 (
            .O(N__47352),
            .I(N__46979));
    SRMux I__11171 (
            .O(N__47351),
            .I(N__46979));
    SRMux I__11170 (
            .O(N__47350),
            .I(N__46979));
    SRMux I__11169 (
            .O(N__47349),
            .I(N__46979));
    SRMux I__11168 (
            .O(N__47348),
            .I(N__46979));
    SRMux I__11167 (
            .O(N__47347),
            .I(N__46979));
    SRMux I__11166 (
            .O(N__47346),
            .I(N__46979));
    SRMux I__11165 (
            .O(N__47345),
            .I(N__46979));
    SRMux I__11164 (
            .O(N__47344),
            .I(N__46979));
    SRMux I__11163 (
            .O(N__47343),
            .I(N__46979));
    SRMux I__11162 (
            .O(N__47342),
            .I(N__46979));
    SRMux I__11161 (
            .O(N__47341),
            .I(N__46979));
    SRMux I__11160 (
            .O(N__47340),
            .I(N__46979));
    SRMux I__11159 (
            .O(N__47339),
            .I(N__46979));
    SRMux I__11158 (
            .O(N__47338),
            .I(N__46979));
    SRMux I__11157 (
            .O(N__47337),
            .I(N__46979));
    SRMux I__11156 (
            .O(N__47336),
            .I(N__46979));
    SRMux I__11155 (
            .O(N__47335),
            .I(N__46979));
    Glb2LocalMux I__11154 (
            .O(N__47332),
            .I(N__46979));
    SRMux I__11153 (
            .O(N__47331),
            .I(N__46979));
    SRMux I__11152 (
            .O(N__47330),
            .I(N__46979));
    SRMux I__11151 (
            .O(N__47329),
            .I(N__46979));
    SRMux I__11150 (
            .O(N__47328),
            .I(N__46979));
    SRMux I__11149 (
            .O(N__47327),
            .I(N__46979));
    SRMux I__11148 (
            .O(N__47326),
            .I(N__46979));
    SRMux I__11147 (
            .O(N__47325),
            .I(N__46979));
    SRMux I__11146 (
            .O(N__47324),
            .I(N__46979));
    SRMux I__11145 (
            .O(N__47323),
            .I(N__46979));
    SRMux I__11144 (
            .O(N__47322),
            .I(N__46979));
    SRMux I__11143 (
            .O(N__47321),
            .I(N__46979));
    SRMux I__11142 (
            .O(N__47320),
            .I(N__46979));
    SRMux I__11141 (
            .O(N__47319),
            .I(N__46979));
    SRMux I__11140 (
            .O(N__47318),
            .I(N__46979));
    SRMux I__11139 (
            .O(N__47317),
            .I(N__46979));
    SRMux I__11138 (
            .O(N__47316),
            .I(N__46979));
    SRMux I__11137 (
            .O(N__47315),
            .I(N__46979));
    SRMux I__11136 (
            .O(N__47314),
            .I(N__46979));
    SRMux I__11135 (
            .O(N__47313),
            .I(N__46979));
    SRMux I__11134 (
            .O(N__47312),
            .I(N__46979));
    SRMux I__11133 (
            .O(N__47311),
            .I(N__46979));
    SRMux I__11132 (
            .O(N__47310),
            .I(N__46979));
    SRMux I__11131 (
            .O(N__47309),
            .I(N__46979));
    SRMux I__11130 (
            .O(N__47308),
            .I(N__46979));
    SRMux I__11129 (
            .O(N__47307),
            .I(N__46979));
    SRMux I__11128 (
            .O(N__47306),
            .I(N__46979));
    SRMux I__11127 (
            .O(N__47305),
            .I(N__46979));
    SRMux I__11126 (
            .O(N__47304),
            .I(N__46979));
    SRMux I__11125 (
            .O(N__47303),
            .I(N__46979));
    SRMux I__11124 (
            .O(N__47302),
            .I(N__46979));
    SRMux I__11123 (
            .O(N__47301),
            .I(N__46979));
    SRMux I__11122 (
            .O(N__47300),
            .I(N__46979));
    SRMux I__11121 (
            .O(N__47299),
            .I(N__46979));
    SRMux I__11120 (
            .O(N__47298),
            .I(N__46979));
    SRMux I__11119 (
            .O(N__47297),
            .I(N__46979));
    SRMux I__11118 (
            .O(N__47296),
            .I(N__46979));
    SRMux I__11117 (
            .O(N__47295),
            .I(N__46979));
    SRMux I__11116 (
            .O(N__47294),
            .I(N__46979));
    SRMux I__11115 (
            .O(N__47293),
            .I(N__46979));
    SRMux I__11114 (
            .O(N__47292),
            .I(N__46979));
    SRMux I__11113 (
            .O(N__47291),
            .I(N__46979));
    SRMux I__11112 (
            .O(N__47290),
            .I(N__46979));
    SRMux I__11111 (
            .O(N__47289),
            .I(N__46979));
    SRMux I__11110 (
            .O(N__47288),
            .I(N__46979));
    SRMux I__11109 (
            .O(N__47287),
            .I(N__46979));
    SRMux I__11108 (
            .O(N__47286),
            .I(N__46979));
    Glb2LocalMux I__11107 (
            .O(N__47283),
            .I(N__46979));
    Glb2LocalMux I__11106 (
            .O(N__47280),
            .I(N__46979));
    SRMux I__11105 (
            .O(N__47279),
            .I(N__46979));
    SRMux I__11104 (
            .O(N__47278),
            .I(N__46979));
    SRMux I__11103 (
            .O(N__47277),
            .I(N__46979));
    SRMux I__11102 (
            .O(N__47276),
            .I(N__46979));
    SRMux I__11101 (
            .O(N__47275),
            .I(N__46979));
    SRMux I__11100 (
            .O(N__47274),
            .I(N__46979));
    SRMux I__11099 (
            .O(N__47273),
            .I(N__46979));
    SRMux I__11098 (
            .O(N__47272),
            .I(N__46979));
    GlobalMux I__11097 (
            .O(N__46979),
            .I(N__46976));
    gio2CtrlBuf I__11096 (
            .O(N__46976),
            .I(red_c_g));
    CascadeMux I__11095 (
            .O(N__46973),
            .I(N__46970));
    InMux I__11094 (
            .O(N__46970),
            .I(N__46966));
    InMux I__11093 (
            .O(N__46969),
            .I(N__46963));
    LocalMux I__11092 (
            .O(N__46966),
            .I(N__46960));
    LocalMux I__11091 (
            .O(N__46963),
            .I(N__46957));
    Span4Mux_h I__11090 (
            .O(N__46960),
            .I(N__46954));
    Span4Mux_h I__11089 (
            .O(N__46957),
            .I(N__46951));
    Odrv4 I__11088 (
            .O(N__46954),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    Odrv4 I__11087 (
            .O(N__46951),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__11086 (
            .O(N__46946),
            .I(N__46942));
    InMux I__11085 (
            .O(N__46945),
            .I(N__46938));
    LocalMux I__11084 (
            .O(N__46942),
            .I(N__46935));
    InMux I__11083 (
            .O(N__46941),
            .I(N__46932));
    LocalMux I__11082 (
            .O(N__46938),
            .I(N__46929));
    Span4Mux_v I__11081 (
            .O(N__46935),
            .I(N__46924));
    LocalMux I__11080 (
            .O(N__46932),
            .I(N__46924));
    Span4Mux_h I__11079 (
            .O(N__46929),
            .I(N__46919));
    Span4Mux_h I__11078 (
            .O(N__46924),
            .I(N__46919));
    Odrv4 I__11077 (
            .O(N__46919),
            .I(measured_delay_tr_5));
    InMux I__11076 (
            .O(N__46916),
            .I(N__46911));
    InMux I__11075 (
            .O(N__46915),
            .I(N__46906));
    InMux I__11074 (
            .O(N__46914),
            .I(N__46906));
    LocalMux I__11073 (
            .O(N__46911),
            .I(N__46903));
    LocalMux I__11072 (
            .O(N__46906),
            .I(N__46900));
    Span4Mux_v I__11071 (
            .O(N__46903),
            .I(N__46897));
    Span4Mux_h I__11070 (
            .O(N__46900),
            .I(N__46894));
    Odrv4 I__11069 (
            .O(N__46897),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    Odrv4 I__11068 (
            .O(N__46894),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    CascadeMux I__11067 (
            .O(N__46889),
            .I(N__46885));
    CascadeMux I__11066 (
            .O(N__46888),
            .I(N__46881));
    InMux I__11065 (
            .O(N__46885),
            .I(N__46878));
    InMux I__11064 (
            .O(N__46884),
            .I(N__46875));
    InMux I__11063 (
            .O(N__46881),
            .I(N__46872));
    LocalMux I__11062 (
            .O(N__46878),
            .I(N__46867));
    LocalMux I__11061 (
            .O(N__46875),
            .I(N__46867));
    LocalMux I__11060 (
            .O(N__46872),
            .I(N__46864));
    Span4Mux_h I__11059 (
            .O(N__46867),
            .I(N__46861));
    Span4Mux_h I__11058 (
            .O(N__46864),
            .I(N__46858));
    Span4Mux_v I__11057 (
            .O(N__46861),
            .I(N__46855));
    Odrv4 I__11056 (
            .O(N__46858),
            .I(measured_delay_tr_3));
    Odrv4 I__11055 (
            .O(N__46855),
            .I(measured_delay_tr_3));
    CascadeMux I__11054 (
            .O(N__46850),
            .I(N__46846));
    InMux I__11053 (
            .O(N__46849),
            .I(N__46843));
    InMux I__11052 (
            .O(N__46846),
            .I(N__46840));
    LocalMux I__11051 (
            .O(N__46843),
            .I(N__46837));
    LocalMux I__11050 (
            .O(N__46840),
            .I(N__46834));
    Span4Mux_h I__11049 (
            .O(N__46837),
            .I(N__46831));
    Span4Mux_h I__11048 (
            .O(N__46834),
            .I(N__46828));
    Odrv4 I__11047 (
            .O(N__46831),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    Odrv4 I__11046 (
            .O(N__46828),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__11045 (
            .O(N__46823),
            .I(N__46819));
    InMux I__11044 (
            .O(N__46822),
            .I(N__46816));
    LocalMux I__11043 (
            .O(N__46819),
            .I(N__46812));
    LocalMux I__11042 (
            .O(N__46816),
            .I(N__46809));
    InMux I__11041 (
            .O(N__46815),
            .I(N__46806));
    Span4Mux_v I__11040 (
            .O(N__46812),
            .I(N__46803));
    Span4Mux_v I__11039 (
            .O(N__46809),
            .I(N__46798));
    LocalMux I__11038 (
            .O(N__46806),
            .I(N__46798));
    Span4Mux_h I__11037 (
            .O(N__46803),
            .I(N__46795));
    Span4Mux_h I__11036 (
            .O(N__46798),
            .I(N__46792));
    Odrv4 I__11035 (
            .O(N__46795),
            .I(measured_delay_tr_8));
    Odrv4 I__11034 (
            .O(N__46792),
            .I(measured_delay_tr_8));
    InMux I__11033 (
            .O(N__46787),
            .I(N__46783));
    InMux I__11032 (
            .O(N__46786),
            .I(N__46780));
    LocalMux I__11031 (
            .O(N__46783),
            .I(N__46777));
    LocalMux I__11030 (
            .O(N__46780),
            .I(N__46774));
    Span4Mux_v I__11029 (
            .O(N__46777),
            .I(N__46771));
    Span4Mux_h I__11028 (
            .O(N__46774),
            .I(N__46768));
    Odrv4 I__11027 (
            .O(N__46771),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv4 I__11026 (
            .O(N__46768),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__11025 (
            .O(N__46763),
            .I(N__46760));
    LocalMux I__11024 (
            .O(N__46760),
            .I(N__46755));
    InMux I__11023 (
            .O(N__46759),
            .I(N__46752));
    InMux I__11022 (
            .O(N__46758),
            .I(N__46749));
    Span4Mux_v I__11021 (
            .O(N__46755),
            .I(N__46742));
    LocalMux I__11020 (
            .O(N__46752),
            .I(N__46742));
    LocalMux I__11019 (
            .O(N__46749),
            .I(N__46742));
    Span4Mux_h I__11018 (
            .O(N__46742),
            .I(N__46739));
    Odrv4 I__11017 (
            .O(N__46739),
            .I(measured_delay_tr_7));
    InMux I__11016 (
            .O(N__46736),
            .I(N__46731));
    InMux I__11015 (
            .O(N__46735),
            .I(N__46728));
    CascadeMux I__11014 (
            .O(N__46734),
            .I(N__46725));
    LocalMux I__11013 (
            .O(N__46731),
            .I(N__46722));
    LocalMux I__11012 (
            .O(N__46728),
            .I(N__46719));
    InMux I__11011 (
            .O(N__46725),
            .I(N__46716));
    Span4Mux_h I__11010 (
            .O(N__46722),
            .I(N__46713));
    Span4Mux_h I__11009 (
            .O(N__46719),
            .I(N__46710));
    LocalMux I__11008 (
            .O(N__46716),
            .I(N__46707));
    Odrv4 I__11007 (
            .O(N__46713),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__11006 (
            .O(N__46710),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv12 I__11005 (
            .O(N__46707),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__11004 (
            .O(N__46700),
            .I(N__46696));
    CascadeMux I__11003 (
            .O(N__46699),
            .I(N__46693));
    LocalMux I__11002 (
            .O(N__46696),
            .I(N__46690));
    InMux I__11001 (
            .O(N__46693),
            .I(N__46687));
    Span4Mux_v I__11000 (
            .O(N__46690),
            .I(N__46682));
    LocalMux I__10999 (
            .O(N__46687),
            .I(N__46682));
    Odrv4 I__10998 (
            .O(N__46682),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__10997 (
            .O(N__46679),
            .I(N__46675));
    CascadeMux I__10996 (
            .O(N__46678),
            .I(N__46671));
    LocalMux I__10995 (
            .O(N__46675),
            .I(N__46668));
    InMux I__10994 (
            .O(N__46674),
            .I(N__46665));
    InMux I__10993 (
            .O(N__46671),
            .I(N__46662));
    Span4Mux_v I__10992 (
            .O(N__46668),
            .I(N__46655));
    LocalMux I__10991 (
            .O(N__46665),
            .I(N__46655));
    LocalMux I__10990 (
            .O(N__46662),
            .I(N__46655));
    Span4Mux_v I__10989 (
            .O(N__46655),
            .I(N__46652));
    Odrv4 I__10988 (
            .O(N__46652),
            .I(measured_delay_tr_13));
    InMux I__10987 (
            .O(N__46649),
            .I(N__46644));
    InMux I__10986 (
            .O(N__46648),
            .I(N__46641));
    InMux I__10985 (
            .O(N__46647),
            .I(N__46638));
    LocalMux I__10984 (
            .O(N__46644),
            .I(N__46630));
    LocalMux I__10983 (
            .O(N__46641),
            .I(N__46630));
    LocalMux I__10982 (
            .O(N__46638),
            .I(N__46630));
    InMux I__10981 (
            .O(N__46637),
            .I(N__46627));
    Span4Mux_v I__10980 (
            .O(N__46630),
            .I(N__46622));
    LocalMux I__10979 (
            .O(N__46627),
            .I(N__46622));
    Odrv4 I__10978 (
            .O(N__46622),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    InMux I__10977 (
            .O(N__46619),
            .I(N__46616));
    LocalMux I__10976 (
            .O(N__46616),
            .I(N__46611));
    InMux I__10975 (
            .O(N__46615),
            .I(N__46608));
    InMux I__10974 (
            .O(N__46614),
            .I(N__46605));
    Span4Mux_v I__10973 (
            .O(N__46611),
            .I(N__46598));
    LocalMux I__10972 (
            .O(N__46608),
            .I(N__46598));
    LocalMux I__10971 (
            .O(N__46605),
            .I(N__46598));
    Span4Mux_h I__10970 (
            .O(N__46598),
            .I(N__46595));
    Odrv4 I__10969 (
            .O(N__46595),
            .I(measured_delay_tr_6));
    InMux I__10968 (
            .O(N__46592),
            .I(N__46588));
    InMux I__10967 (
            .O(N__46591),
            .I(N__46585));
    LocalMux I__10966 (
            .O(N__46588),
            .I(N__46582));
    LocalMux I__10965 (
            .O(N__46585),
            .I(N__46579));
    Span4Mux_v I__10964 (
            .O(N__46582),
            .I(N__46576));
    Span4Mux_h I__10963 (
            .O(N__46579),
            .I(N__46573));
    Odrv4 I__10962 (
            .O(N__46576),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    Odrv4 I__10961 (
            .O(N__46573),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__10960 (
            .O(N__46568),
            .I(N__46565));
    LocalMux I__10959 (
            .O(N__46565),
            .I(N__46560));
    InMux I__10958 (
            .O(N__46564),
            .I(N__46557));
    InMux I__10957 (
            .O(N__46563),
            .I(N__46554));
    Span4Mux_v I__10956 (
            .O(N__46560),
            .I(N__46547));
    LocalMux I__10955 (
            .O(N__46557),
            .I(N__46547));
    LocalMux I__10954 (
            .O(N__46554),
            .I(N__46547));
    Span4Mux_h I__10953 (
            .O(N__46547),
            .I(N__46544));
    Odrv4 I__10952 (
            .O(N__46544),
            .I(measured_delay_tr_4));
    InMux I__10951 (
            .O(N__46541),
            .I(N__46525));
    InMux I__10950 (
            .O(N__46540),
            .I(N__46525));
    InMux I__10949 (
            .O(N__46539),
            .I(N__46525));
    InMux I__10948 (
            .O(N__46538),
            .I(N__46525));
    InMux I__10947 (
            .O(N__46537),
            .I(N__46516));
    InMux I__10946 (
            .O(N__46536),
            .I(N__46516));
    InMux I__10945 (
            .O(N__46535),
            .I(N__46516));
    InMux I__10944 (
            .O(N__46534),
            .I(N__46516));
    LocalMux I__10943 (
            .O(N__46525),
            .I(N__46513));
    LocalMux I__10942 (
            .O(N__46516),
            .I(N__46510));
    Span4Mux_h I__10941 (
            .O(N__46513),
            .I(N__46507));
    Span4Mux_h I__10940 (
            .O(N__46510),
            .I(N__46504));
    Odrv4 I__10939 (
            .O(N__46507),
            .I(\delay_measurement_inst.N_324 ));
    Odrv4 I__10938 (
            .O(N__46504),
            .I(\delay_measurement_inst.N_324 ));
    InMux I__10937 (
            .O(N__46499),
            .I(N__46490));
    InMux I__10936 (
            .O(N__46498),
            .I(N__46490));
    InMux I__10935 (
            .O(N__46497),
            .I(N__46490));
    LocalMux I__10934 (
            .O(N__46490),
            .I(N__46484));
    InMux I__10933 (
            .O(N__46489),
            .I(N__46477));
    InMux I__10932 (
            .O(N__46488),
            .I(N__46477));
    InMux I__10931 (
            .O(N__46487),
            .I(N__46477));
    Odrv4 I__10930 (
            .O(N__46484),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6 ));
    LocalMux I__10929 (
            .O(N__46477),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6 ));
    InMux I__10928 (
            .O(N__46472),
            .I(N__46469));
    LocalMux I__10927 (
            .O(N__46469),
            .I(N__46464));
    CascadeMux I__10926 (
            .O(N__46468),
            .I(N__46461));
    InMux I__10925 (
            .O(N__46467),
            .I(N__46458));
    Span4Mux_h I__10924 (
            .O(N__46464),
            .I(N__46455));
    InMux I__10923 (
            .O(N__46461),
            .I(N__46452));
    LocalMux I__10922 (
            .O(N__46458),
            .I(N__46449));
    Span4Mux_v I__10921 (
            .O(N__46455),
            .I(N__46444));
    LocalMux I__10920 (
            .O(N__46452),
            .I(N__46444));
    Span4Mux_h I__10919 (
            .O(N__46449),
            .I(N__46441));
    Span4Mux_h I__10918 (
            .O(N__46444),
            .I(N__46438));
    Odrv4 I__10917 (
            .O(N__46441),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__10916 (
            .O(N__46438),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    CascadeMux I__10915 (
            .O(N__46433),
            .I(N__46429));
    CascadeMux I__10914 (
            .O(N__46432),
            .I(N__46426));
    InMux I__10913 (
            .O(N__46429),
            .I(N__46423));
    InMux I__10912 (
            .O(N__46426),
            .I(N__46419));
    LocalMux I__10911 (
            .O(N__46423),
            .I(N__46416));
    InMux I__10910 (
            .O(N__46422),
            .I(N__46413));
    LocalMux I__10909 (
            .O(N__46419),
            .I(N__46410));
    Span4Mux_h I__10908 (
            .O(N__46416),
            .I(N__46405));
    LocalMux I__10907 (
            .O(N__46413),
            .I(N__46405));
    Span4Mux_h I__10906 (
            .O(N__46410),
            .I(N__46402));
    Span4Mux_v I__10905 (
            .O(N__46405),
            .I(N__46399));
    Odrv4 I__10904 (
            .O(N__46402),
            .I(measured_delay_tr_2));
    Odrv4 I__10903 (
            .O(N__46399),
            .I(measured_delay_tr_2));
    CascadeMux I__10902 (
            .O(N__46394),
            .I(\delay_measurement_inst.delay_tr_timer.N_331_cascade_ ));
    InMux I__10901 (
            .O(N__46391),
            .I(N__46388));
    LocalMux I__10900 (
            .O(N__46388),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ));
    InMux I__10899 (
            .O(N__46385),
            .I(N__46382));
    LocalMux I__10898 (
            .O(N__46382),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ));
    CascadeMux I__10897 (
            .O(N__46379),
            .I(\delay_measurement_inst.delay_tr_timer.N_321_cascade_ ));
    InMux I__10896 (
            .O(N__46376),
            .I(N__46372));
    InMux I__10895 (
            .O(N__46375),
            .I(N__46369));
    LocalMux I__10894 (
            .O(N__46372),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14 ));
    LocalMux I__10893 (
            .O(N__46369),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14 ));
    InMux I__10892 (
            .O(N__46364),
            .I(N__46358));
    InMux I__10891 (
            .O(N__46363),
            .I(N__46358));
    LocalMux I__10890 (
            .O(N__46358),
            .I(\delay_measurement_inst.delay_tr_timer.N_331 ));
    InMux I__10889 (
            .O(N__46355),
            .I(N__46352));
    LocalMux I__10888 (
            .O(N__46352),
            .I(\delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14 ));
    InMux I__10887 (
            .O(N__46349),
            .I(N__46345));
    InMux I__10886 (
            .O(N__46348),
            .I(N__46342));
    LocalMux I__10885 (
            .O(N__46345),
            .I(N__46337));
    LocalMux I__10884 (
            .O(N__46342),
            .I(N__46334));
    InMux I__10883 (
            .O(N__46341),
            .I(N__46329));
    InMux I__10882 (
            .O(N__46340),
            .I(N__46329));
    Span4Mux_v I__10881 (
            .O(N__46337),
            .I(N__46322));
    Span4Mux_v I__10880 (
            .O(N__46334),
            .I(N__46322));
    LocalMux I__10879 (
            .O(N__46329),
            .I(N__46322));
    Odrv4 I__10878 (
            .O(N__46322),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    InMux I__10877 (
            .O(N__46319),
            .I(N__46314));
    InMux I__10876 (
            .O(N__46318),
            .I(N__46309));
    InMux I__10875 (
            .O(N__46317),
            .I(N__46306));
    LocalMux I__10874 (
            .O(N__46314),
            .I(N__46303));
    InMux I__10873 (
            .O(N__46313),
            .I(N__46298));
    InMux I__10872 (
            .O(N__46312),
            .I(N__46298));
    LocalMux I__10871 (
            .O(N__46309),
            .I(N__46295));
    LocalMux I__10870 (
            .O(N__46306),
            .I(N__46288));
    Span4Mux_v I__10869 (
            .O(N__46303),
            .I(N__46288));
    LocalMux I__10868 (
            .O(N__46298),
            .I(N__46288));
    Span12Mux_v I__10867 (
            .O(N__46295),
            .I(N__46285));
    Span4Mux_v I__10866 (
            .O(N__46288),
            .I(N__46282));
    Odrv12 I__10865 (
            .O(N__46285),
            .I(measured_delay_tr_14));
    Odrv4 I__10864 (
            .O(N__46282),
            .I(measured_delay_tr_14));
    InMux I__10863 (
            .O(N__46277),
            .I(N__46269));
    CascadeMux I__10862 (
            .O(N__46276),
            .I(N__46266));
    InMux I__10861 (
            .O(N__46275),
            .I(N__46263));
    InMux I__10860 (
            .O(N__46274),
            .I(N__46260));
    InMux I__10859 (
            .O(N__46273),
            .I(N__46255));
    InMux I__10858 (
            .O(N__46272),
            .I(N__46255));
    LocalMux I__10857 (
            .O(N__46269),
            .I(N__46251));
    InMux I__10856 (
            .O(N__46266),
            .I(N__46248));
    LocalMux I__10855 (
            .O(N__46263),
            .I(N__46241));
    LocalMux I__10854 (
            .O(N__46260),
            .I(N__46241));
    LocalMux I__10853 (
            .O(N__46255),
            .I(N__46241));
    InMux I__10852 (
            .O(N__46254),
            .I(N__46238));
    Span4Mux_v I__10851 (
            .O(N__46251),
            .I(N__46235));
    LocalMux I__10850 (
            .O(N__46248),
            .I(N__46232));
    Span4Mux_v I__10849 (
            .O(N__46241),
            .I(N__46229));
    LocalMux I__10848 (
            .O(N__46238),
            .I(N__46226));
    Odrv4 I__10847 (
            .O(N__46235),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv4 I__10846 (
            .O(N__46232),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv4 I__10845 (
            .O(N__46229),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv12 I__10844 (
            .O(N__46226),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    CascadeMux I__10843 (
            .O(N__46217),
            .I(N__46214));
    InMux I__10842 (
            .O(N__46214),
            .I(N__46210));
    InMux I__10841 (
            .O(N__46213),
            .I(N__46207));
    LocalMux I__10840 (
            .O(N__46210),
            .I(N__46201));
    LocalMux I__10839 (
            .O(N__46207),
            .I(N__46198));
    InMux I__10838 (
            .O(N__46206),
            .I(N__46191));
    InMux I__10837 (
            .O(N__46205),
            .I(N__46191));
    InMux I__10836 (
            .O(N__46204),
            .I(N__46191));
    Odrv4 I__10835 (
            .O(N__46201),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ));
    Odrv12 I__10834 (
            .O(N__46198),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ));
    LocalMux I__10833 (
            .O(N__46191),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ));
    CascadeMux I__10832 (
            .O(N__46184),
            .I(N__46174));
    InMux I__10831 (
            .O(N__46183),
            .I(N__46170));
    InMux I__10830 (
            .O(N__46182),
            .I(N__46167));
    InMux I__10829 (
            .O(N__46181),
            .I(N__46164));
    InMux I__10828 (
            .O(N__46180),
            .I(N__46161));
    InMux I__10827 (
            .O(N__46179),
            .I(N__46156));
    InMux I__10826 (
            .O(N__46178),
            .I(N__46156));
    CascadeMux I__10825 (
            .O(N__46177),
            .I(N__46152));
    InMux I__10824 (
            .O(N__46174),
            .I(N__46149));
    InMux I__10823 (
            .O(N__46173),
            .I(N__46146));
    LocalMux I__10822 (
            .O(N__46170),
            .I(N__46143));
    LocalMux I__10821 (
            .O(N__46167),
            .I(N__46140));
    LocalMux I__10820 (
            .O(N__46164),
            .I(N__46137));
    LocalMux I__10819 (
            .O(N__46161),
            .I(N__46132));
    LocalMux I__10818 (
            .O(N__46156),
            .I(N__46132));
    InMux I__10817 (
            .O(N__46155),
            .I(N__46127));
    InMux I__10816 (
            .O(N__46152),
            .I(N__46127));
    LocalMux I__10815 (
            .O(N__46149),
            .I(N__46120));
    LocalMux I__10814 (
            .O(N__46146),
            .I(N__46120));
    Span4Mux_v I__10813 (
            .O(N__46143),
            .I(N__46120));
    Span4Mux_v I__10812 (
            .O(N__46140),
            .I(N__46115));
    Span4Mux_v I__10811 (
            .O(N__46137),
            .I(N__46115));
    Span4Mux_v I__10810 (
            .O(N__46132),
            .I(N__46110));
    LocalMux I__10809 (
            .O(N__46127),
            .I(N__46110));
    Span4Mux_h I__10808 (
            .O(N__46120),
            .I(N__46105));
    Span4Mux_h I__10807 (
            .O(N__46115),
            .I(N__46105));
    Span4Mux_v I__10806 (
            .O(N__46110),
            .I(N__46102));
    Span4Mux_v I__10805 (
            .O(N__46105),
            .I(N__46099));
    Span4Mux_h I__10804 (
            .O(N__46102),
            .I(N__46096));
    Odrv4 I__10803 (
            .O(N__46099),
            .I(measured_delay_tr_15));
    Odrv4 I__10802 (
            .O(N__46096),
            .I(measured_delay_tr_15));
    InMux I__10801 (
            .O(N__46091),
            .I(N__46087));
    InMux I__10800 (
            .O(N__46090),
            .I(N__46084));
    LocalMux I__10799 (
            .O(N__46087),
            .I(N__46081));
    LocalMux I__10798 (
            .O(N__46084),
            .I(N__46078));
    Span4Mux_v I__10797 (
            .O(N__46081),
            .I(N__46075));
    Span4Mux_h I__10796 (
            .O(N__46078),
            .I(N__46072));
    Odrv4 I__10795 (
            .O(N__46075),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    Odrv4 I__10794 (
            .O(N__46072),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    CascadeMux I__10793 (
            .O(N__46067),
            .I(N__46064));
    InMux I__10792 (
            .O(N__46064),
            .I(N__46061));
    LocalMux I__10791 (
            .O(N__46061),
            .I(N__46057));
    CascadeMux I__10790 (
            .O(N__46060),
            .I(N__46054));
    Span4Mux_v I__10789 (
            .O(N__46057),
            .I(N__46051));
    InMux I__10788 (
            .O(N__46054),
            .I(N__46048));
    Span4Mux_h I__10787 (
            .O(N__46051),
            .I(N__46043));
    LocalMux I__10786 (
            .O(N__46048),
            .I(N__46043));
    Span4Mux_h I__10785 (
            .O(N__46043),
            .I(N__46040));
    Odrv4 I__10784 (
            .O(N__46040),
            .I(measured_delay_tr_1));
    CascadeMux I__10783 (
            .O(N__46037),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ));
    InMux I__10782 (
            .O(N__46034),
            .I(N__46031));
    LocalMux I__10781 (
            .O(N__46031),
            .I(N__46025));
    InMux I__10780 (
            .O(N__46030),
            .I(N__46022));
    InMux I__10779 (
            .O(N__46029),
            .I(N__46018));
    InMux I__10778 (
            .O(N__46028),
            .I(N__46015));
    Span4Mux_v I__10777 (
            .O(N__46025),
            .I(N__46012));
    LocalMux I__10776 (
            .O(N__46022),
            .I(N__46009));
    InMux I__10775 (
            .O(N__46021),
            .I(N__46006));
    LocalMux I__10774 (
            .O(N__46018),
            .I(N__46003));
    LocalMux I__10773 (
            .O(N__46015),
            .I(N__46000));
    Span4Mux_v I__10772 (
            .O(N__46012),
            .I(N__45993));
    Span4Mux_v I__10771 (
            .O(N__46009),
            .I(N__45993));
    LocalMux I__10770 (
            .O(N__46006),
            .I(N__45993));
    Odrv4 I__10769 (
            .O(N__46003),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__10768 (
            .O(N__46000),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__10767 (
            .O(N__45993),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    CascadeMux I__10766 (
            .O(N__45986),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_ ));
    InMux I__10765 (
            .O(N__45983),
            .I(N__45980));
    LocalMux I__10764 (
            .O(N__45980),
            .I(\delay_measurement_inst.delay_tr_timer.N_320_4 ));
    CascadeMux I__10763 (
            .O(N__45977),
            .I(\delay_measurement_inst.delay_tr_timer.N_320_4_cascade_ ));
    InMux I__10762 (
            .O(N__45974),
            .I(N__45971));
    LocalMux I__10761 (
            .O(N__45971),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ));
    InMux I__10760 (
            .O(N__45968),
            .I(N__45965));
    LocalMux I__10759 (
            .O(N__45965),
            .I(N__45961));
    InMux I__10758 (
            .O(N__45964),
            .I(N__45958));
    Span4Mux_v I__10757 (
            .O(N__45961),
            .I(N__45953));
    LocalMux I__10756 (
            .O(N__45958),
            .I(N__45953));
    Odrv4 I__10755 (
            .O(N__45953),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__10754 (
            .O(N__45950),
            .I(N__45946));
    InMux I__10753 (
            .O(N__45949),
            .I(N__45943));
    LocalMux I__10752 (
            .O(N__45946),
            .I(N__45940));
    LocalMux I__10751 (
            .O(N__45943),
            .I(N__45937));
    Span4Mux_v I__10750 (
            .O(N__45940),
            .I(N__45934));
    Span4Mux_h I__10749 (
            .O(N__45937),
            .I(N__45931));
    Odrv4 I__10748 (
            .O(N__45934),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    Odrv4 I__10747 (
            .O(N__45931),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__10746 (
            .O(N__45926),
            .I(N__45922));
    InMux I__10745 (
            .O(N__45925),
            .I(N__45919));
    LocalMux I__10744 (
            .O(N__45922),
            .I(N__45916));
    LocalMux I__10743 (
            .O(N__45919),
            .I(N__45913));
    Span4Mux_h I__10742 (
            .O(N__45916),
            .I(N__45909));
    Span4Mux_h I__10741 (
            .O(N__45913),
            .I(N__45906));
    InMux I__10740 (
            .O(N__45912),
            .I(N__45903));
    Odrv4 I__10739 (
            .O(N__45909),
            .I(\delay_measurement_inst.N_328 ));
    Odrv4 I__10738 (
            .O(N__45906),
            .I(\delay_measurement_inst.N_328 ));
    LocalMux I__10737 (
            .O(N__45903),
            .I(\delay_measurement_inst.N_328 ));
    InMux I__10736 (
            .O(N__45896),
            .I(N__45893));
    LocalMux I__10735 (
            .O(N__45893),
            .I(N__45890));
    Span4Mux_h I__10734 (
            .O(N__45890),
            .I(N__45886));
    InMux I__10733 (
            .O(N__45889),
            .I(N__45883));
    Odrv4 I__10732 (
            .O(N__45886),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__10731 (
            .O(N__45883),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__10730 (
            .O(N__45878),
            .I(N__45875));
    LocalMux I__10729 (
            .O(N__45875),
            .I(N__45872));
    Span4Mux_v I__10728 (
            .O(N__45872),
            .I(N__45869));
    Odrv4 I__10727 (
            .O(N__45869),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__10726 (
            .O(N__45866),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__10725 (
            .O(N__45863),
            .I(N__45860));
    LocalMux I__10724 (
            .O(N__45860),
            .I(N__45856));
    InMux I__10723 (
            .O(N__45859),
            .I(N__45853));
    Span4Mux_h I__10722 (
            .O(N__45856),
            .I(N__45850));
    LocalMux I__10721 (
            .O(N__45853),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__10720 (
            .O(N__45850),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__10719 (
            .O(N__45845),
            .I(N__45842));
    LocalMux I__10718 (
            .O(N__45842),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__10717 (
            .O(N__45839),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__10716 (
            .O(N__45836),
            .I(N__45833));
    LocalMux I__10715 (
            .O(N__45833),
            .I(N__45829));
    InMux I__10714 (
            .O(N__45832),
            .I(N__45826));
    Span4Mux_v I__10713 (
            .O(N__45829),
            .I(N__45823));
    LocalMux I__10712 (
            .O(N__45826),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__10711 (
            .O(N__45823),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__10710 (
            .O(N__45818),
            .I(N__45815));
    LocalMux I__10709 (
            .O(N__45815),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__10708 (
            .O(N__45812),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__10707 (
            .O(N__45809),
            .I(N__45806));
    LocalMux I__10706 (
            .O(N__45806),
            .I(N__45802));
    InMux I__10705 (
            .O(N__45805),
            .I(N__45799));
    Span4Mux_h I__10704 (
            .O(N__45802),
            .I(N__45796));
    LocalMux I__10703 (
            .O(N__45799),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__10702 (
            .O(N__45796),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__10701 (
            .O(N__45791),
            .I(N__45788));
    LocalMux I__10700 (
            .O(N__45788),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__10699 (
            .O(N__45785),
            .I(bfn_18_21_0_));
    InMux I__10698 (
            .O(N__45782),
            .I(N__45779));
    LocalMux I__10697 (
            .O(N__45779),
            .I(N__45775));
    InMux I__10696 (
            .O(N__45778),
            .I(N__45772));
    Span4Mux_h I__10695 (
            .O(N__45775),
            .I(N__45769));
    LocalMux I__10694 (
            .O(N__45772),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__10693 (
            .O(N__45769),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__10692 (
            .O(N__45764),
            .I(N__45761));
    LocalMux I__10691 (
            .O(N__45761),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__10690 (
            .O(N__45758),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__10689 (
            .O(N__45755),
            .I(N__45752));
    LocalMux I__10688 (
            .O(N__45752),
            .I(N__45748));
    InMux I__10687 (
            .O(N__45751),
            .I(N__45745));
    Span4Mux_h I__10686 (
            .O(N__45748),
            .I(N__45742));
    LocalMux I__10685 (
            .O(N__45745),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__10684 (
            .O(N__45742),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__10683 (
            .O(N__45737),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__10682 (
            .O(N__45734),
            .I(N__45731));
    LocalMux I__10681 (
            .O(N__45731),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__10680 (
            .O(N__45728),
            .I(N__45725));
    LocalMux I__10679 (
            .O(N__45725),
            .I(N__45721));
    InMux I__10678 (
            .O(N__45724),
            .I(N__45718));
    Odrv4 I__10677 (
            .O(N__45721),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ));
    LocalMux I__10676 (
            .O(N__45718),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ));
    InMux I__10675 (
            .O(N__45713),
            .I(N__45709));
    InMux I__10674 (
            .O(N__45712),
            .I(N__45705));
    LocalMux I__10673 (
            .O(N__45709),
            .I(N__45702));
    InMux I__10672 (
            .O(N__45708),
            .I(N__45699));
    LocalMux I__10671 (
            .O(N__45705),
            .I(N__45696));
    Span4Mux_h I__10670 (
            .O(N__45702),
            .I(N__45686));
    LocalMux I__10669 (
            .O(N__45699),
            .I(N__45686));
    Span4Mux_h I__10668 (
            .O(N__45696),
            .I(N__45686));
    InMux I__10667 (
            .O(N__45695),
            .I(N__45683));
    InMux I__10666 (
            .O(N__45694),
            .I(N__45680));
    InMux I__10665 (
            .O(N__45693),
            .I(N__45677));
    Odrv4 I__10664 (
            .O(N__45686),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    LocalMux I__10663 (
            .O(N__45683),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    LocalMux I__10662 (
            .O(N__45680),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    LocalMux I__10661 (
            .O(N__45677),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    CascadeMux I__10660 (
            .O(N__45668),
            .I(N__45665));
    InMux I__10659 (
            .O(N__45665),
            .I(N__45662));
    LocalMux I__10658 (
            .O(N__45662),
            .I(N__45659));
    Span4Mux_h I__10657 (
            .O(N__45659),
            .I(N__45656));
    Odrv4 I__10656 (
            .O(N__45656),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__10655 (
            .O(N__45653),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__10654 (
            .O(N__45650),
            .I(N__45647));
    LocalMux I__10653 (
            .O(N__45647),
            .I(N__45644));
    Span4Mux_v I__10652 (
            .O(N__45644),
            .I(N__45640));
    InMux I__10651 (
            .O(N__45643),
            .I(N__45637));
    Odrv4 I__10650 (
            .O(N__45640),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__10649 (
            .O(N__45637),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__10648 (
            .O(N__45632),
            .I(N__45629));
    LocalMux I__10647 (
            .O(N__45629),
            .I(N__45626));
    Span4Mux_h I__10646 (
            .O(N__45626),
            .I(N__45623));
    Odrv4 I__10645 (
            .O(N__45623),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__10644 (
            .O(N__45620),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__10643 (
            .O(N__45617),
            .I(N__45614));
    LocalMux I__10642 (
            .O(N__45614),
            .I(N__45611));
    Span4Mux_h I__10641 (
            .O(N__45611),
            .I(N__45607));
    InMux I__10640 (
            .O(N__45610),
            .I(N__45604));
    Odrv4 I__10639 (
            .O(N__45607),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__10638 (
            .O(N__45604),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__10637 (
            .O(N__45599),
            .I(N__45596));
    InMux I__10636 (
            .O(N__45596),
            .I(N__45593));
    LocalMux I__10635 (
            .O(N__45593),
            .I(N__45590));
    Span4Mux_h I__10634 (
            .O(N__45590),
            .I(N__45587));
    Odrv4 I__10633 (
            .O(N__45587),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__10632 (
            .O(N__45584),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__10631 (
            .O(N__45581),
            .I(N__45578));
    LocalMux I__10630 (
            .O(N__45578),
            .I(N__45574));
    InMux I__10629 (
            .O(N__45577),
            .I(N__45571));
    Span4Mux_h I__10628 (
            .O(N__45574),
            .I(N__45568));
    LocalMux I__10627 (
            .O(N__45571),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__10626 (
            .O(N__45568),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__10625 (
            .O(N__45563),
            .I(N__45560));
    LocalMux I__10624 (
            .O(N__45560),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__10623 (
            .O(N__45557),
            .I(bfn_18_20_0_));
    InMux I__10622 (
            .O(N__45554),
            .I(N__45551));
    LocalMux I__10621 (
            .O(N__45551),
            .I(N__45548));
    Span4Mux_h I__10620 (
            .O(N__45548),
            .I(N__45544));
    InMux I__10619 (
            .O(N__45547),
            .I(N__45541));
    Odrv4 I__10618 (
            .O(N__45544),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__10617 (
            .O(N__45541),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__10616 (
            .O(N__45536),
            .I(N__45533));
    InMux I__10615 (
            .O(N__45533),
            .I(N__45530));
    LocalMux I__10614 (
            .O(N__45530),
            .I(N__45527));
    Span4Mux_h I__10613 (
            .O(N__45527),
            .I(N__45524));
    Odrv4 I__10612 (
            .O(N__45524),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__10611 (
            .O(N__45521),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__10610 (
            .O(N__45518),
            .I(N__45515));
    LocalMux I__10609 (
            .O(N__45515),
            .I(N__45511));
    InMux I__10608 (
            .O(N__45514),
            .I(N__45508));
    Span4Mux_h I__10607 (
            .O(N__45511),
            .I(N__45505));
    LocalMux I__10606 (
            .O(N__45508),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__10605 (
            .O(N__45505),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__10604 (
            .O(N__45500),
            .I(N__45497));
    LocalMux I__10603 (
            .O(N__45497),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__10602 (
            .O(N__45494),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__10601 (
            .O(N__45491),
            .I(N__45488));
    LocalMux I__10600 (
            .O(N__45488),
            .I(N__45484));
    InMux I__10599 (
            .O(N__45487),
            .I(N__45481));
    Span4Mux_h I__10598 (
            .O(N__45484),
            .I(N__45478));
    LocalMux I__10597 (
            .O(N__45481),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__10596 (
            .O(N__45478),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__10595 (
            .O(N__45473),
            .I(N__45470));
    LocalMux I__10594 (
            .O(N__45470),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__10593 (
            .O(N__45467),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__10592 (
            .O(N__45464),
            .I(N__45461));
    LocalMux I__10591 (
            .O(N__45461),
            .I(N__45457));
    InMux I__10590 (
            .O(N__45460),
            .I(N__45454));
    Span4Mux_v I__10589 (
            .O(N__45457),
            .I(N__45451));
    LocalMux I__10588 (
            .O(N__45454),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__10587 (
            .O(N__45451),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__10586 (
            .O(N__45446),
            .I(N__45443));
    LocalMux I__10585 (
            .O(N__45443),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__10584 (
            .O(N__45440),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__10583 (
            .O(N__45437),
            .I(N__45430));
    InMux I__10582 (
            .O(N__45436),
            .I(N__45430));
    InMux I__10581 (
            .O(N__45435),
            .I(N__45427));
    LocalMux I__10580 (
            .O(N__45430),
            .I(N__45424));
    LocalMux I__10579 (
            .O(N__45427),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__10578 (
            .O(N__45424),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    CascadeMux I__10577 (
            .O(N__45419),
            .I(N__45416));
    InMux I__10576 (
            .O(N__45416),
            .I(N__45412));
    InMux I__10575 (
            .O(N__45415),
            .I(N__45409));
    LocalMux I__10574 (
            .O(N__45412),
            .I(N__45406));
    LocalMux I__10573 (
            .O(N__45409),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__10572 (
            .O(N__45406),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    InMux I__10571 (
            .O(N__45401),
            .I(N__45398));
    LocalMux I__10570 (
            .O(N__45398),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__10569 (
            .O(N__45395),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__10568 (
            .O(N__45392),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__10567 (
            .O(N__45389),
            .I(N__45384));
    CEMux I__10566 (
            .O(N__45388),
            .I(N__45381));
    CEMux I__10565 (
            .O(N__45387),
            .I(N__45378));
    LocalMux I__10564 (
            .O(N__45384),
            .I(N__45374));
    LocalMux I__10563 (
            .O(N__45381),
            .I(N__45370));
    LocalMux I__10562 (
            .O(N__45378),
            .I(N__45367));
    CEMux I__10561 (
            .O(N__45377),
            .I(N__45364));
    Span4Mux_v I__10560 (
            .O(N__45374),
            .I(N__45361));
    CEMux I__10559 (
            .O(N__45373),
            .I(N__45358));
    Span4Mux_v I__10558 (
            .O(N__45370),
            .I(N__45347));
    Span4Mux_v I__10557 (
            .O(N__45367),
            .I(N__45347));
    LocalMux I__10556 (
            .O(N__45364),
            .I(N__45347));
    Span4Mux_v I__10555 (
            .O(N__45361),
            .I(N__45347));
    LocalMux I__10554 (
            .O(N__45358),
            .I(N__45347));
    Span4Mux_v I__10553 (
            .O(N__45347),
            .I(N__45344));
    Span4Mux_h I__10552 (
            .O(N__45344),
            .I(N__45341));
    Odrv4 I__10551 (
            .O(N__45341),
            .I(\delay_measurement_inst.delay_tr_timer.N_337_i ));
    InMux I__10550 (
            .O(N__45338),
            .I(N__45335));
    LocalMux I__10549 (
            .O(N__45335),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__10548 (
            .O(N__45332),
            .I(N__45329));
    InMux I__10547 (
            .O(N__45329),
            .I(N__45324));
    InMux I__10546 (
            .O(N__45328),
            .I(N__45321));
    InMux I__10545 (
            .O(N__45327),
            .I(N__45318));
    LocalMux I__10544 (
            .O(N__45324),
            .I(N__45315));
    LocalMux I__10543 (
            .O(N__45321),
            .I(N__45310));
    LocalMux I__10542 (
            .O(N__45318),
            .I(N__45310));
    Span4Mux_h I__10541 (
            .O(N__45315),
            .I(N__45305));
    Span4Mux_v I__10540 (
            .O(N__45310),
            .I(N__45305));
    Odrv4 I__10539 (
            .O(N__45305),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__10538 (
            .O(N__45302),
            .I(N__45299));
    LocalMux I__10537 (
            .O(N__45299),
            .I(N__45296));
    Span4Mux_h I__10536 (
            .O(N__45296),
            .I(N__45292));
    InMux I__10535 (
            .O(N__45295),
            .I(N__45289));
    Odrv4 I__10534 (
            .O(N__45292),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__10533 (
            .O(N__45289),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__10532 (
            .O(N__45284),
            .I(N__45281));
    LocalMux I__10531 (
            .O(N__45281),
            .I(N__45278));
    Span4Mux_h I__10530 (
            .O(N__45278),
            .I(N__45275));
    Odrv4 I__10529 (
            .O(N__45275),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__10528 (
            .O(N__45272),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__10527 (
            .O(N__45269),
            .I(N__45266));
    LocalMux I__10526 (
            .O(N__45266),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ));
    CascadeMux I__10525 (
            .O(N__45263),
            .I(N__45260));
    InMux I__10524 (
            .O(N__45260),
            .I(N__45257));
    LocalMux I__10523 (
            .O(N__45257),
            .I(N__45254));
    Span4Mux_v I__10522 (
            .O(N__45254),
            .I(N__45250));
    InMux I__10521 (
            .O(N__45253),
            .I(N__45247));
    Odrv4 I__10520 (
            .O(N__45250),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__10519 (
            .O(N__45247),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__10518 (
            .O(N__45242),
            .I(N__45239));
    LocalMux I__10517 (
            .O(N__45239),
            .I(N__45236));
    Span12Mux_h I__10516 (
            .O(N__45236),
            .I(N__45233));
    Odrv12 I__10515 (
            .O(N__45233),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__10514 (
            .O(N__45230),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__10513 (
            .O(N__45227),
            .I(N__45224));
    LocalMux I__10512 (
            .O(N__45224),
            .I(N__45221));
    Span4Mux_h I__10511 (
            .O(N__45221),
            .I(N__45217));
    InMux I__10510 (
            .O(N__45220),
            .I(N__45214));
    Odrv4 I__10509 (
            .O(N__45217),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__10508 (
            .O(N__45214),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__10507 (
            .O(N__45209),
            .I(N__45206));
    LocalMux I__10506 (
            .O(N__45206),
            .I(N__45203));
    Span4Mux_v I__10505 (
            .O(N__45203),
            .I(N__45200));
    Odrv4 I__10504 (
            .O(N__45200),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__10503 (
            .O(N__45197),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__10502 (
            .O(N__45194),
            .I(N__45191));
    LocalMux I__10501 (
            .O(N__45191),
            .I(N__45188));
    Span4Mux_v I__10500 (
            .O(N__45188),
            .I(N__45184));
    InMux I__10499 (
            .O(N__45187),
            .I(N__45181));
    Odrv4 I__10498 (
            .O(N__45184),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__10497 (
            .O(N__45181),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__10496 (
            .O(N__45176),
            .I(N__45173));
    InMux I__10495 (
            .O(N__45173),
            .I(N__45170));
    LocalMux I__10494 (
            .O(N__45170),
            .I(N__45167));
    Span4Mux_h I__10493 (
            .O(N__45167),
            .I(N__45164));
    Odrv4 I__10492 (
            .O(N__45164),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__10491 (
            .O(N__45161),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__10490 (
            .O(N__45158),
            .I(N__45155));
    LocalMux I__10489 (
            .O(N__45155),
            .I(N__45152));
    Span4Mux_h I__10488 (
            .O(N__45152),
            .I(N__45148));
    InMux I__10487 (
            .O(N__45151),
            .I(N__45145));
    Odrv4 I__10486 (
            .O(N__45148),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__10485 (
            .O(N__45145),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__10484 (
            .O(N__45140),
            .I(N__45136));
    CascadeMux I__10483 (
            .O(N__45139),
            .I(N__45133));
    InMux I__10482 (
            .O(N__45136),
            .I(N__45127));
    InMux I__10481 (
            .O(N__45133),
            .I(N__45127));
    InMux I__10480 (
            .O(N__45132),
            .I(N__45124));
    LocalMux I__10479 (
            .O(N__45127),
            .I(N__45121));
    LocalMux I__10478 (
            .O(N__45124),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__10477 (
            .O(N__45121),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__10476 (
            .O(N__45116),
            .I(N__45113));
    LocalMux I__10475 (
            .O(N__45113),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__10474 (
            .O(N__45110),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__10473 (
            .O(N__45107),
            .I(N__45101));
    InMux I__10472 (
            .O(N__45106),
            .I(N__45101));
    LocalMux I__10471 (
            .O(N__45101),
            .I(N__45097));
    InMux I__10470 (
            .O(N__45100),
            .I(N__45094));
    Span4Mux_h I__10469 (
            .O(N__45097),
            .I(N__45091));
    LocalMux I__10468 (
            .O(N__45094),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__10467 (
            .O(N__45091),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__10466 (
            .O(N__45086),
            .I(N__45083));
    LocalMux I__10465 (
            .O(N__45083),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__10464 (
            .O(N__45080),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__10463 (
            .O(N__45077),
            .I(N__45074));
    InMux I__10462 (
            .O(N__45074),
            .I(N__45070));
    InMux I__10461 (
            .O(N__45073),
            .I(N__45067));
    LocalMux I__10460 (
            .O(N__45070),
            .I(N__45061));
    LocalMux I__10459 (
            .O(N__45067),
            .I(N__45061));
    InMux I__10458 (
            .O(N__45066),
            .I(N__45058));
    Span4Mux_v I__10457 (
            .O(N__45061),
            .I(N__45055));
    LocalMux I__10456 (
            .O(N__45058),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__10455 (
            .O(N__45055),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    CascadeMux I__10454 (
            .O(N__45050),
            .I(N__45047));
    InMux I__10453 (
            .O(N__45047),
            .I(N__45044));
    LocalMux I__10452 (
            .O(N__45044),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__10451 (
            .O(N__45041),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__10450 (
            .O(N__45038),
            .I(N__45034));
    InMux I__10449 (
            .O(N__45037),
            .I(N__45031));
    InMux I__10448 (
            .O(N__45034),
            .I(N__45028));
    LocalMux I__10447 (
            .O(N__45031),
            .I(N__45022));
    LocalMux I__10446 (
            .O(N__45028),
            .I(N__45022));
    InMux I__10445 (
            .O(N__45027),
            .I(N__45019));
    Span4Mux_v I__10444 (
            .O(N__45022),
            .I(N__45016));
    LocalMux I__10443 (
            .O(N__45019),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__10442 (
            .O(N__45016),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__10441 (
            .O(N__45011),
            .I(N__45008));
    LocalMux I__10440 (
            .O(N__45008),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__10439 (
            .O(N__45005),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__10438 (
            .O(N__45002),
            .I(N__44995));
    InMux I__10437 (
            .O(N__45001),
            .I(N__44995));
    InMux I__10436 (
            .O(N__45000),
            .I(N__44992));
    LocalMux I__10435 (
            .O(N__44995),
            .I(N__44989));
    LocalMux I__10434 (
            .O(N__44992),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__10433 (
            .O(N__44989),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__10432 (
            .O(N__44984),
            .I(N__44981));
    LocalMux I__10431 (
            .O(N__44981),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__10430 (
            .O(N__44978),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__10429 (
            .O(N__44975),
            .I(N__44972));
    LocalMux I__10428 (
            .O(N__44972),
            .I(N__44968));
    CascadeMux I__10427 (
            .O(N__44971),
            .I(N__44964));
    Span4Mux_h I__10426 (
            .O(N__44968),
            .I(N__44961));
    InMux I__10425 (
            .O(N__44967),
            .I(N__44958));
    InMux I__10424 (
            .O(N__44964),
            .I(N__44955));
    Odrv4 I__10423 (
            .O(N__44961),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__10422 (
            .O(N__44958),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__10421 (
            .O(N__44955),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__10420 (
            .O(N__44948),
            .I(N__44945));
    LocalMux I__10419 (
            .O(N__44945),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__10418 (
            .O(N__44942),
            .I(bfn_18_18_0_));
    CascadeMux I__10417 (
            .O(N__44939),
            .I(N__44936));
    InMux I__10416 (
            .O(N__44936),
            .I(N__44933));
    LocalMux I__10415 (
            .O(N__44933),
            .I(N__44928));
    CascadeMux I__10414 (
            .O(N__44932),
            .I(N__44925));
    InMux I__10413 (
            .O(N__44931),
            .I(N__44922));
    Span4Mux_h I__10412 (
            .O(N__44928),
            .I(N__44919));
    InMux I__10411 (
            .O(N__44925),
            .I(N__44916));
    LocalMux I__10410 (
            .O(N__44922),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__10409 (
            .O(N__44919),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__10408 (
            .O(N__44916),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    CascadeMux I__10407 (
            .O(N__44909),
            .I(N__44906));
    InMux I__10406 (
            .O(N__44906),
            .I(N__44903));
    LocalMux I__10405 (
            .O(N__44903),
            .I(N__44900));
    Odrv4 I__10404 (
            .O(N__44900),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10403 (
            .O(N__44897),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__10402 (
            .O(N__44894),
            .I(N__44890));
    InMux I__10401 (
            .O(N__44893),
            .I(N__44887));
    LocalMux I__10400 (
            .O(N__44890),
            .I(N__44884));
    LocalMux I__10399 (
            .O(N__44887),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__10398 (
            .O(N__44884),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__10397 (
            .O(N__44879),
            .I(N__44875));
    CascadeMux I__10396 (
            .O(N__44878),
            .I(N__44872));
    InMux I__10395 (
            .O(N__44875),
            .I(N__44866));
    InMux I__10394 (
            .O(N__44872),
            .I(N__44866));
    InMux I__10393 (
            .O(N__44871),
            .I(N__44863));
    LocalMux I__10392 (
            .O(N__44866),
            .I(N__44860));
    LocalMux I__10391 (
            .O(N__44863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__10390 (
            .O(N__44860),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__10389 (
            .O(N__44855),
            .I(N__44852));
    LocalMux I__10388 (
            .O(N__44852),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__10387 (
            .O(N__44849),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__10386 (
            .O(N__44846),
            .I(N__44842));
    InMux I__10385 (
            .O(N__44845),
            .I(N__44839));
    InMux I__10384 (
            .O(N__44842),
            .I(N__44836));
    LocalMux I__10383 (
            .O(N__44839),
            .I(N__44830));
    LocalMux I__10382 (
            .O(N__44836),
            .I(N__44830));
    InMux I__10381 (
            .O(N__44835),
            .I(N__44827));
    Span4Mux_v I__10380 (
            .O(N__44830),
            .I(N__44824));
    LocalMux I__10379 (
            .O(N__44827),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__10378 (
            .O(N__44824),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__10377 (
            .O(N__44819),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__10376 (
            .O(N__44816),
            .I(N__44812));
    CascadeMux I__10375 (
            .O(N__44815),
            .I(N__44809));
    InMux I__10374 (
            .O(N__44812),
            .I(N__44803));
    InMux I__10373 (
            .O(N__44809),
            .I(N__44803));
    InMux I__10372 (
            .O(N__44808),
            .I(N__44800));
    LocalMux I__10371 (
            .O(N__44803),
            .I(N__44797));
    LocalMux I__10370 (
            .O(N__44800),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__10369 (
            .O(N__44797),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__10368 (
            .O(N__44792),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__10367 (
            .O(N__44789),
            .I(N__44785));
    CascadeMux I__10366 (
            .O(N__44788),
            .I(N__44782));
    InMux I__10365 (
            .O(N__44785),
            .I(N__44776));
    InMux I__10364 (
            .O(N__44782),
            .I(N__44776));
    InMux I__10363 (
            .O(N__44781),
            .I(N__44773));
    LocalMux I__10362 (
            .O(N__44776),
            .I(N__44770));
    LocalMux I__10361 (
            .O(N__44773),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__10360 (
            .O(N__44770),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__10359 (
            .O(N__44765),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__10358 (
            .O(N__44762),
            .I(N__44755));
    InMux I__10357 (
            .O(N__44761),
            .I(N__44755));
    InMux I__10356 (
            .O(N__44760),
            .I(N__44752));
    LocalMux I__10355 (
            .O(N__44755),
            .I(N__44749));
    LocalMux I__10354 (
            .O(N__44752),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__10353 (
            .O(N__44749),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__10352 (
            .O(N__44744),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__10351 (
            .O(N__44741),
            .I(N__44734));
    InMux I__10350 (
            .O(N__44740),
            .I(N__44734));
    InMux I__10349 (
            .O(N__44739),
            .I(N__44731));
    LocalMux I__10348 (
            .O(N__44734),
            .I(N__44728));
    LocalMux I__10347 (
            .O(N__44731),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__10346 (
            .O(N__44728),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__10345 (
            .O(N__44723),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__10344 (
            .O(N__44720),
            .I(N__44716));
    InMux I__10343 (
            .O(N__44719),
            .I(N__44712));
    InMux I__10342 (
            .O(N__44716),
            .I(N__44709));
    InMux I__10341 (
            .O(N__44715),
            .I(N__44706));
    LocalMux I__10340 (
            .O(N__44712),
            .I(N__44701));
    LocalMux I__10339 (
            .O(N__44709),
            .I(N__44701));
    LocalMux I__10338 (
            .O(N__44706),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__10337 (
            .O(N__44701),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__10336 (
            .O(N__44696),
            .I(bfn_18_17_0_));
    InMux I__10335 (
            .O(N__44693),
            .I(N__44689));
    CascadeMux I__10334 (
            .O(N__44692),
            .I(N__44685));
    LocalMux I__10333 (
            .O(N__44689),
            .I(N__44682));
    InMux I__10332 (
            .O(N__44688),
            .I(N__44679));
    InMux I__10331 (
            .O(N__44685),
            .I(N__44676));
    Odrv4 I__10330 (
            .O(N__44682),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__10329 (
            .O(N__44679),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__10328 (
            .O(N__44676),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__10327 (
            .O(N__44669),
            .I(N__44666));
    LocalMux I__10326 (
            .O(N__44666),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__10325 (
            .O(N__44663),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__10324 (
            .O(N__44660),
            .I(N__44656));
    CascadeMux I__10323 (
            .O(N__44659),
            .I(N__44653));
    InMux I__10322 (
            .O(N__44656),
            .I(N__44647));
    InMux I__10321 (
            .O(N__44653),
            .I(N__44647));
    InMux I__10320 (
            .O(N__44652),
            .I(N__44644));
    LocalMux I__10319 (
            .O(N__44647),
            .I(N__44641));
    LocalMux I__10318 (
            .O(N__44644),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__10317 (
            .O(N__44641),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__10316 (
            .O(N__44636),
            .I(N__44633));
    LocalMux I__10315 (
            .O(N__44633),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__10314 (
            .O(N__44630),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__10313 (
            .O(N__44627),
            .I(N__44623));
    CascadeMux I__10312 (
            .O(N__44626),
            .I(N__44620));
    InMux I__10311 (
            .O(N__44623),
            .I(N__44614));
    InMux I__10310 (
            .O(N__44620),
            .I(N__44614));
    InMux I__10309 (
            .O(N__44619),
            .I(N__44611));
    LocalMux I__10308 (
            .O(N__44614),
            .I(N__44608));
    LocalMux I__10307 (
            .O(N__44611),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__10306 (
            .O(N__44608),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__10305 (
            .O(N__44603),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__10304 (
            .O(N__44600),
            .I(N__44596));
    CascadeMux I__10303 (
            .O(N__44599),
            .I(N__44593));
    InMux I__10302 (
            .O(N__44596),
            .I(N__44587));
    InMux I__10301 (
            .O(N__44593),
            .I(N__44587));
    InMux I__10300 (
            .O(N__44592),
            .I(N__44584));
    LocalMux I__10299 (
            .O(N__44587),
            .I(N__44581));
    LocalMux I__10298 (
            .O(N__44584),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__10297 (
            .O(N__44581),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__10296 (
            .O(N__44576),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__10295 (
            .O(N__44573),
            .I(N__44567));
    InMux I__10294 (
            .O(N__44572),
            .I(N__44567));
    LocalMux I__10293 (
            .O(N__44567),
            .I(N__44563));
    InMux I__10292 (
            .O(N__44566),
            .I(N__44560));
    Span4Mux_h I__10291 (
            .O(N__44563),
            .I(N__44557));
    LocalMux I__10290 (
            .O(N__44560),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__10289 (
            .O(N__44557),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__10288 (
            .O(N__44552),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__10287 (
            .O(N__44549),
            .I(N__44543));
    InMux I__10286 (
            .O(N__44548),
            .I(N__44543));
    LocalMux I__10285 (
            .O(N__44543),
            .I(N__44539));
    InMux I__10284 (
            .O(N__44542),
            .I(N__44536));
    Span4Mux_h I__10283 (
            .O(N__44539),
            .I(N__44533));
    LocalMux I__10282 (
            .O(N__44536),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__10281 (
            .O(N__44533),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__10280 (
            .O(N__44528),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__10279 (
            .O(N__44525),
            .I(N__44521));
    InMux I__10278 (
            .O(N__44524),
            .I(N__44518));
    InMux I__10277 (
            .O(N__44521),
            .I(N__44515));
    LocalMux I__10276 (
            .O(N__44518),
            .I(N__44509));
    LocalMux I__10275 (
            .O(N__44515),
            .I(N__44509));
    InMux I__10274 (
            .O(N__44514),
            .I(N__44506));
    Span4Mux_v I__10273 (
            .O(N__44509),
            .I(N__44503));
    LocalMux I__10272 (
            .O(N__44506),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__10271 (
            .O(N__44503),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__10270 (
            .O(N__44498),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__10269 (
            .O(N__44495),
            .I(N__44491));
    CascadeMux I__10268 (
            .O(N__44494),
            .I(N__44488));
    InMux I__10267 (
            .O(N__44491),
            .I(N__44483));
    InMux I__10266 (
            .O(N__44488),
            .I(N__44483));
    LocalMux I__10265 (
            .O(N__44483),
            .I(N__44479));
    InMux I__10264 (
            .O(N__44482),
            .I(N__44476));
    Span4Mux_v I__10263 (
            .O(N__44479),
            .I(N__44473));
    LocalMux I__10262 (
            .O(N__44476),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__10261 (
            .O(N__44473),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__10260 (
            .O(N__44468),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__10259 (
            .O(N__44465),
            .I(N__44462));
    LocalMux I__10258 (
            .O(N__44462),
            .I(N__44458));
    CascadeMux I__10257 (
            .O(N__44461),
            .I(N__44454));
    Span4Mux_h I__10256 (
            .O(N__44458),
            .I(N__44451));
    InMux I__10255 (
            .O(N__44457),
            .I(N__44448));
    InMux I__10254 (
            .O(N__44454),
            .I(N__44445));
    Odrv4 I__10253 (
            .O(N__44451),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__10252 (
            .O(N__44448),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__10251 (
            .O(N__44445),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__10250 (
            .O(N__44438),
            .I(bfn_18_16_0_));
    InMux I__10249 (
            .O(N__44435),
            .I(N__44432));
    LocalMux I__10248 (
            .O(N__44432),
            .I(N__44427));
    InMux I__10247 (
            .O(N__44431),
            .I(N__44424));
    InMux I__10246 (
            .O(N__44430),
            .I(N__44421));
    Odrv4 I__10245 (
            .O(N__44427),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__10244 (
            .O(N__44424),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__10243 (
            .O(N__44421),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__10242 (
            .O(N__44414),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10241 (
            .O(N__44411),
            .I(N__44407));
    InMux I__10240 (
            .O(N__44410),
            .I(N__44404));
    InMux I__10239 (
            .O(N__44407),
            .I(N__44401));
    LocalMux I__10238 (
            .O(N__44404),
            .I(N__44395));
    LocalMux I__10237 (
            .O(N__44401),
            .I(N__44395));
    InMux I__10236 (
            .O(N__44400),
            .I(N__44392));
    Span4Mux_v I__10235 (
            .O(N__44395),
            .I(N__44389));
    LocalMux I__10234 (
            .O(N__44392),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__10233 (
            .O(N__44389),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__10232 (
            .O(N__44384),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__10231 (
            .O(N__44381),
            .I(N__44378));
    LocalMux I__10230 (
            .O(N__44378),
            .I(N__44375));
    Span4Mux_h I__10229 (
            .O(N__44375),
            .I(N__44370));
    InMux I__10228 (
            .O(N__44374),
            .I(N__44367));
    InMux I__10227 (
            .O(N__44373),
            .I(N__44364));
    Odrv4 I__10226 (
            .O(N__44370),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__10225 (
            .O(N__44367),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__10224 (
            .O(N__44364),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__10223 (
            .O(N__44357),
            .I(N__44352));
    InMux I__10222 (
            .O(N__44356),
            .I(N__44349));
    InMux I__10221 (
            .O(N__44355),
            .I(N__44346));
    LocalMux I__10220 (
            .O(N__44352),
            .I(N__44341));
    LocalMux I__10219 (
            .O(N__44349),
            .I(N__44341));
    LocalMux I__10218 (
            .O(N__44346),
            .I(N__44336));
    Span4Mux_v I__10217 (
            .O(N__44341),
            .I(N__44336));
    Odrv4 I__10216 (
            .O(N__44336),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    CEMux I__10215 (
            .O(N__44333),
            .I(N__44315));
    CEMux I__10214 (
            .O(N__44332),
            .I(N__44315));
    CEMux I__10213 (
            .O(N__44331),
            .I(N__44315));
    CEMux I__10212 (
            .O(N__44330),
            .I(N__44315));
    CEMux I__10211 (
            .O(N__44329),
            .I(N__44315));
    CEMux I__10210 (
            .O(N__44328),
            .I(N__44315));
    GlobalMux I__10209 (
            .O(N__44315),
            .I(N__44312));
    gio2CtrlBuf I__10208 (
            .O(N__44312),
            .I(\delay_measurement_inst.delay_hc_timer.N_335_i_g ));
    InMux I__10207 (
            .O(N__44309),
            .I(N__44306));
    LocalMux I__10206 (
            .O(N__44306),
            .I(N__44302));
    InMux I__10205 (
            .O(N__44305),
            .I(N__44299));
    Span4Mux_v I__10204 (
            .O(N__44302),
            .I(N__44293));
    LocalMux I__10203 (
            .O(N__44299),
            .I(N__44293));
    InMux I__10202 (
            .O(N__44298),
            .I(N__44290));
    Odrv4 I__10201 (
            .O(N__44293),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__10200 (
            .O(N__44290),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__10199 (
            .O(N__44285),
            .I(N__44281));
    InMux I__10198 (
            .O(N__44284),
            .I(N__44278));
    LocalMux I__10197 (
            .O(N__44281),
            .I(N__44274));
    LocalMux I__10196 (
            .O(N__44278),
            .I(N__44271));
    InMux I__10195 (
            .O(N__44277),
            .I(N__44268));
    Odrv12 I__10194 (
            .O(N__44274),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    Odrv4 I__10193 (
            .O(N__44271),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__10192 (
            .O(N__44268),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    CascadeMux I__10191 (
            .O(N__44261),
            .I(N__44258));
    InMux I__10190 (
            .O(N__44258),
            .I(N__44254));
    InMux I__10189 (
            .O(N__44257),
            .I(N__44251));
    LocalMux I__10188 (
            .O(N__44254),
            .I(N__44247));
    LocalMux I__10187 (
            .O(N__44251),
            .I(N__44244));
    CascadeMux I__10186 (
            .O(N__44250),
            .I(N__44241));
    Span4Mux_v I__10185 (
            .O(N__44247),
            .I(N__44236));
    Span4Mux_v I__10184 (
            .O(N__44244),
            .I(N__44236));
    InMux I__10183 (
            .O(N__44241),
            .I(N__44233));
    Odrv4 I__10182 (
            .O(N__44236),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    LocalMux I__10181 (
            .O(N__44233),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__10180 (
            .O(N__44228),
            .I(N__44224));
    InMux I__10179 (
            .O(N__44227),
            .I(N__44221));
    LocalMux I__10178 (
            .O(N__44224),
            .I(N__44217));
    LocalMux I__10177 (
            .O(N__44221),
            .I(N__44214));
    InMux I__10176 (
            .O(N__44220),
            .I(N__44211));
    Odrv12 I__10175 (
            .O(N__44217),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    Odrv4 I__10174 (
            .O(N__44214),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__10173 (
            .O(N__44211),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__10172 (
            .O(N__44204),
            .I(N__44201));
    LocalMux I__10171 (
            .O(N__44201),
            .I(N__44197));
    InMux I__10170 (
            .O(N__44200),
            .I(N__44194));
    Span4Mux_v I__10169 (
            .O(N__44197),
            .I(N__44189));
    LocalMux I__10168 (
            .O(N__44194),
            .I(N__44189));
    Span4Mux_v I__10167 (
            .O(N__44189),
            .I(N__44186));
    Sp12to4 I__10166 (
            .O(N__44186),
            .I(N__44178));
    InMux I__10165 (
            .O(N__44185),
            .I(N__44175));
    InMux I__10164 (
            .O(N__44184),
            .I(N__44168));
    InMux I__10163 (
            .O(N__44183),
            .I(N__44168));
    InMux I__10162 (
            .O(N__44182),
            .I(N__44168));
    InMux I__10161 (
            .O(N__44181),
            .I(N__44165));
    Odrv12 I__10160 (
            .O(N__44178),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__10159 (
            .O(N__44175),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__10158 (
            .O(N__44168),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__10157 (
            .O(N__44165),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    InMux I__10156 (
            .O(N__44156),
            .I(N__44153));
    LocalMux I__10155 (
            .O(N__44153),
            .I(N__44150));
    Span4Mux_h I__10154 (
            .O(N__44150),
            .I(N__44146));
    InMux I__10153 (
            .O(N__44149),
            .I(N__44142));
    Span4Mux_h I__10152 (
            .O(N__44146),
            .I(N__44139));
    InMux I__10151 (
            .O(N__44145),
            .I(N__44135));
    LocalMux I__10150 (
            .O(N__44142),
            .I(N__44130));
    Span4Mux_v I__10149 (
            .O(N__44139),
            .I(N__44127));
    InMux I__10148 (
            .O(N__44138),
            .I(N__44124));
    LocalMux I__10147 (
            .O(N__44135),
            .I(N__44121));
    InMux I__10146 (
            .O(N__44134),
            .I(N__44118));
    InMux I__10145 (
            .O(N__44133),
            .I(N__44115));
    Span4Mux_h I__10144 (
            .O(N__44130),
            .I(N__44112));
    Span4Mux_v I__10143 (
            .O(N__44127),
            .I(N__44107));
    LocalMux I__10142 (
            .O(N__44124),
            .I(N__44107));
    Span4Mux_v I__10141 (
            .O(N__44121),
            .I(N__44102));
    LocalMux I__10140 (
            .O(N__44118),
            .I(N__44102));
    LocalMux I__10139 (
            .O(N__44115),
            .I(N__44099));
    Odrv4 I__10138 (
            .O(N__44112),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    Odrv4 I__10137 (
            .O(N__44107),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    Odrv4 I__10136 (
            .O(N__44102),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    Odrv4 I__10135 (
            .O(N__44099),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__10134 (
            .O(N__44090),
            .I(N__44087));
    LocalMux I__10133 (
            .O(N__44087),
            .I(N__44084));
    Odrv4 I__10132 (
            .O(N__44084),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1 ));
    InMux I__10131 (
            .O(N__44081),
            .I(N__44075));
    InMux I__10130 (
            .O(N__44080),
            .I(N__44072));
    InMux I__10129 (
            .O(N__44079),
            .I(N__44068));
    InMux I__10128 (
            .O(N__44078),
            .I(N__44064));
    LocalMux I__10127 (
            .O(N__44075),
            .I(N__44061));
    LocalMux I__10126 (
            .O(N__44072),
            .I(N__44058));
    InMux I__10125 (
            .O(N__44071),
            .I(N__44055));
    LocalMux I__10124 (
            .O(N__44068),
            .I(N__44052));
    InMux I__10123 (
            .O(N__44067),
            .I(N__44049));
    LocalMux I__10122 (
            .O(N__44064),
            .I(N__44046));
    Span4Mux_h I__10121 (
            .O(N__44061),
            .I(N__44043));
    Span4Mux_h I__10120 (
            .O(N__44058),
            .I(N__44040));
    LocalMux I__10119 (
            .O(N__44055),
            .I(N__44037));
    Span4Mux_h I__10118 (
            .O(N__44052),
            .I(N__44032));
    LocalMux I__10117 (
            .O(N__44049),
            .I(N__44032));
    Odrv4 I__10116 (
            .O(N__44046),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__10115 (
            .O(N__44043),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__10114 (
            .O(N__44040),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__10113 (
            .O(N__44037),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__10112 (
            .O(N__44032),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    CascadeMux I__10111 (
            .O(N__44021),
            .I(N__44017));
    InMux I__10110 (
            .O(N__44020),
            .I(N__44010));
    InMux I__10109 (
            .O(N__44017),
            .I(N__44007));
    InMux I__10108 (
            .O(N__44016),
            .I(N__44000));
    InMux I__10107 (
            .O(N__44015),
            .I(N__44000));
    InMux I__10106 (
            .O(N__44014),
            .I(N__44000));
    InMux I__10105 (
            .O(N__44013),
            .I(N__43997));
    LocalMux I__10104 (
            .O(N__44010),
            .I(N__43994));
    LocalMux I__10103 (
            .O(N__44007),
            .I(N__43991));
    LocalMux I__10102 (
            .O(N__44000),
            .I(N__43988));
    LocalMux I__10101 (
            .O(N__43997),
            .I(N__43985));
    Span4Mux_h I__10100 (
            .O(N__43994),
            .I(N__43982));
    Span4Mux_h I__10099 (
            .O(N__43991),
            .I(N__43977));
    Span4Mux_h I__10098 (
            .O(N__43988),
            .I(N__43977));
    Odrv4 I__10097 (
            .O(N__43985),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    Odrv4 I__10096 (
            .O(N__43982),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    Odrv4 I__10095 (
            .O(N__43977),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    CascadeMux I__10094 (
            .O(N__43970),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1_cascade_ ));
    InMux I__10093 (
            .O(N__43967),
            .I(N__43964));
    LocalMux I__10092 (
            .O(N__43964),
            .I(N__43960));
    InMux I__10091 (
            .O(N__43963),
            .I(N__43957));
    Span4Mux_v I__10090 (
            .O(N__43960),
            .I(N__43951));
    LocalMux I__10089 (
            .O(N__43957),
            .I(N__43951));
    InMux I__10088 (
            .O(N__43956),
            .I(N__43947));
    Span4Mux_v I__10087 (
            .O(N__43951),
            .I(N__43944));
    InMux I__10086 (
            .O(N__43950),
            .I(N__43940));
    LocalMux I__10085 (
            .O(N__43947),
            .I(N__43935));
    Span4Mux_h I__10084 (
            .O(N__43944),
            .I(N__43935));
    InMux I__10083 (
            .O(N__43943),
            .I(N__43932));
    LocalMux I__10082 (
            .O(N__43940),
            .I(N__43929));
    Span4Mux_h I__10081 (
            .O(N__43935),
            .I(N__43925));
    LocalMux I__10080 (
            .O(N__43932),
            .I(N__43922));
    Span4Mux_h I__10079 (
            .O(N__43929),
            .I(N__43919));
    InMux I__10078 (
            .O(N__43928),
            .I(N__43916));
    Odrv4 I__10077 (
            .O(N__43925),
            .I(\delay_measurement_inst.delay_hc_reg3lto19_1 ));
    Odrv4 I__10076 (
            .O(N__43922),
            .I(\delay_measurement_inst.delay_hc_reg3lto19_1 ));
    Odrv4 I__10075 (
            .O(N__43919),
            .I(\delay_measurement_inst.delay_hc_reg3lto19_1 ));
    LocalMux I__10074 (
            .O(N__43916),
            .I(\delay_measurement_inst.delay_hc_reg3lto19_1 ));
    InMux I__10073 (
            .O(N__43907),
            .I(N__43904));
    LocalMux I__10072 (
            .O(N__43904),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_2 ));
    InMux I__10071 (
            .O(N__43901),
            .I(N__43897));
    InMux I__10070 (
            .O(N__43900),
            .I(N__43893));
    LocalMux I__10069 (
            .O(N__43897),
            .I(N__43890));
    InMux I__10068 (
            .O(N__43896),
            .I(N__43887));
    LocalMux I__10067 (
            .O(N__43893),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__10066 (
            .O(N__43890),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__10065 (
            .O(N__43887),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__10064 (
            .O(N__43880),
            .I(N__43876));
    InMux I__10063 (
            .O(N__43879),
            .I(N__43872));
    LocalMux I__10062 (
            .O(N__43876),
            .I(N__43869));
    InMux I__10061 (
            .O(N__43875),
            .I(N__43866));
    LocalMux I__10060 (
            .O(N__43872),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__10059 (
            .O(N__43869),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10058 (
            .O(N__43866),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__10057 (
            .O(N__43859),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__10056 (
            .O(N__43856),
            .I(N__43849));
    CascadeMux I__10055 (
            .O(N__43855),
            .I(N__43846));
    InMux I__10054 (
            .O(N__43854),
            .I(N__43836));
    InMux I__10053 (
            .O(N__43853),
            .I(N__43830));
    InMux I__10052 (
            .O(N__43852),
            .I(N__43819));
    InMux I__10051 (
            .O(N__43849),
            .I(N__43816));
    InMux I__10050 (
            .O(N__43846),
            .I(N__43799));
    InMux I__10049 (
            .O(N__43845),
            .I(N__43799));
    InMux I__10048 (
            .O(N__43844),
            .I(N__43799));
    InMux I__10047 (
            .O(N__43843),
            .I(N__43799));
    InMux I__10046 (
            .O(N__43842),
            .I(N__43799));
    InMux I__10045 (
            .O(N__43841),
            .I(N__43799));
    InMux I__10044 (
            .O(N__43840),
            .I(N__43799));
    InMux I__10043 (
            .O(N__43839),
            .I(N__43799));
    LocalMux I__10042 (
            .O(N__43836),
            .I(N__43796));
    InMux I__10041 (
            .O(N__43835),
            .I(N__43791));
    InMux I__10040 (
            .O(N__43834),
            .I(N__43791));
    CascadeMux I__10039 (
            .O(N__43833),
            .I(N__43787));
    LocalMux I__10038 (
            .O(N__43830),
            .I(N__43784));
    InMux I__10037 (
            .O(N__43829),
            .I(N__43767));
    InMux I__10036 (
            .O(N__43828),
            .I(N__43767));
    InMux I__10035 (
            .O(N__43827),
            .I(N__43767));
    InMux I__10034 (
            .O(N__43826),
            .I(N__43767));
    InMux I__10033 (
            .O(N__43825),
            .I(N__43767));
    InMux I__10032 (
            .O(N__43824),
            .I(N__43767));
    InMux I__10031 (
            .O(N__43823),
            .I(N__43767));
    InMux I__10030 (
            .O(N__43822),
            .I(N__43767));
    LocalMux I__10029 (
            .O(N__43819),
            .I(N__43764));
    LocalMux I__10028 (
            .O(N__43816),
            .I(N__43755));
    LocalMux I__10027 (
            .O(N__43799),
            .I(N__43755));
    Span4Mux_v I__10026 (
            .O(N__43796),
            .I(N__43755));
    LocalMux I__10025 (
            .O(N__43791),
            .I(N__43755));
    InMux I__10024 (
            .O(N__43790),
            .I(N__43750));
    InMux I__10023 (
            .O(N__43787),
            .I(N__43750));
    Span4Mux_v I__10022 (
            .O(N__43784),
            .I(N__43747));
    LocalMux I__10021 (
            .O(N__43767),
            .I(N__43740));
    Span4Mux_v I__10020 (
            .O(N__43764),
            .I(N__43740));
    Span4Mux_v I__10019 (
            .O(N__43755),
            .I(N__43740));
    LocalMux I__10018 (
            .O(N__43750),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10017 (
            .O(N__43747),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10016 (
            .O(N__43740),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__10015 (
            .O(N__43733),
            .I(N__43729));
    CascadeMux I__10014 (
            .O(N__43732),
            .I(N__43725));
    InMux I__10013 (
            .O(N__43729),
            .I(N__43715));
    InMux I__10012 (
            .O(N__43728),
            .I(N__43715));
    InMux I__10011 (
            .O(N__43725),
            .I(N__43707));
    CascadeMux I__10010 (
            .O(N__43724),
            .I(N__43704));
    CascadeMux I__10009 (
            .O(N__43723),
            .I(N__43697));
    CascadeMux I__10008 (
            .O(N__43722),
            .I(N__43694));
    CascadeMux I__10007 (
            .O(N__43721),
            .I(N__43691));
    CascadeMux I__10006 (
            .O(N__43720),
            .I(N__43688));
    LocalMux I__10005 (
            .O(N__43715),
            .I(N__43685));
    InMux I__10004 (
            .O(N__43714),
            .I(N__43682));
    CascadeMux I__10003 (
            .O(N__43713),
            .I(N__43678));
    CascadeMux I__10002 (
            .O(N__43712),
            .I(N__43675));
    CascadeMux I__10001 (
            .O(N__43711),
            .I(N__43672));
    CascadeMux I__10000 (
            .O(N__43710),
            .I(N__43669));
    LocalMux I__9999 (
            .O(N__43707),
            .I(N__43661));
    InMux I__9998 (
            .O(N__43704),
            .I(N__43657));
    InMux I__9997 (
            .O(N__43703),
            .I(N__43640));
    InMux I__9996 (
            .O(N__43702),
            .I(N__43640));
    InMux I__9995 (
            .O(N__43701),
            .I(N__43640));
    InMux I__9994 (
            .O(N__43700),
            .I(N__43640));
    InMux I__9993 (
            .O(N__43697),
            .I(N__43640));
    InMux I__9992 (
            .O(N__43694),
            .I(N__43640));
    InMux I__9991 (
            .O(N__43691),
            .I(N__43640));
    InMux I__9990 (
            .O(N__43688),
            .I(N__43640));
    Span4Mux_v I__9989 (
            .O(N__43685),
            .I(N__43635));
    LocalMux I__9988 (
            .O(N__43682),
            .I(N__43635));
    InMux I__9987 (
            .O(N__43681),
            .I(N__43618));
    InMux I__9986 (
            .O(N__43678),
            .I(N__43618));
    InMux I__9985 (
            .O(N__43675),
            .I(N__43618));
    InMux I__9984 (
            .O(N__43672),
            .I(N__43618));
    InMux I__9983 (
            .O(N__43669),
            .I(N__43618));
    InMux I__9982 (
            .O(N__43668),
            .I(N__43618));
    InMux I__9981 (
            .O(N__43667),
            .I(N__43618));
    InMux I__9980 (
            .O(N__43666),
            .I(N__43618));
    InMux I__9979 (
            .O(N__43665),
            .I(N__43613));
    InMux I__9978 (
            .O(N__43664),
            .I(N__43613));
    Span4Mux_v I__9977 (
            .O(N__43661),
            .I(N__43610));
    InMux I__9976 (
            .O(N__43660),
            .I(N__43607));
    LocalMux I__9975 (
            .O(N__43657),
            .I(N__43600));
    LocalMux I__9974 (
            .O(N__43640),
            .I(N__43600));
    Span4Mux_h I__9973 (
            .O(N__43635),
            .I(N__43600));
    LocalMux I__9972 (
            .O(N__43618),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    LocalMux I__9971 (
            .O(N__43613),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9970 (
            .O(N__43610),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    LocalMux I__9969 (
            .O(N__43607),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9968 (
            .O(N__43600),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    CascadeMux I__9967 (
            .O(N__43589),
            .I(N__43580));
    CascadeMux I__9966 (
            .O(N__43588),
            .I(N__43577));
    CascadeMux I__9965 (
            .O(N__43587),
            .I(N__43574));
    CascadeMux I__9964 (
            .O(N__43586),
            .I(N__43565));
    InMux I__9963 (
            .O(N__43585),
            .I(N__43561));
    InMux I__9962 (
            .O(N__43584),
            .I(N__43550));
    InMux I__9961 (
            .O(N__43583),
            .I(N__43547));
    InMux I__9960 (
            .O(N__43580),
            .I(N__43540));
    InMux I__9959 (
            .O(N__43577),
            .I(N__43540));
    InMux I__9958 (
            .O(N__43574),
            .I(N__43540));
    InMux I__9957 (
            .O(N__43573),
            .I(N__43529));
    InMux I__9956 (
            .O(N__43572),
            .I(N__43529));
    InMux I__9955 (
            .O(N__43571),
            .I(N__43529));
    InMux I__9954 (
            .O(N__43570),
            .I(N__43529));
    InMux I__9953 (
            .O(N__43569),
            .I(N__43529));
    InMux I__9952 (
            .O(N__43568),
            .I(N__43526));
    InMux I__9951 (
            .O(N__43565),
            .I(N__43521));
    InMux I__9950 (
            .O(N__43564),
            .I(N__43521));
    LocalMux I__9949 (
            .O(N__43561),
            .I(N__43516));
    InMux I__9948 (
            .O(N__43560),
            .I(N__43499));
    InMux I__9947 (
            .O(N__43559),
            .I(N__43499));
    InMux I__9946 (
            .O(N__43558),
            .I(N__43499));
    InMux I__9945 (
            .O(N__43557),
            .I(N__43499));
    InMux I__9944 (
            .O(N__43556),
            .I(N__43499));
    InMux I__9943 (
            .O(N__43555),
            .I(N__43499));
    InMux I__9942 (
            .O(N__43554),
            .I(N__43499));
    InMux I__9941 (
            .O(N__43553),
            .I(N__43499));
    LocalMux I__9940 (
            .O(N__43550),
            .I(N__43494));
    LocalMux I__9939 (
            .O(N__43547),
            .I(N__43494));
    LocalMux I__9938 (
            .O(N__43540),
            .I(N__43485));
    LocalMux I__9937 (
            .O(N__43529),
            .I(N__43485));
    LocalMux I__9936 (
            .O(N__43526),
            .I(N__43485));
    LocalMux I__9935 (
            .O(N__43521),
            .I(N__43485));
    InMux I__9934 (
            .O(N__43520),
            .I(N__43480));
    InMux I__9933 (
            .O(N__43519),
            .I(N__43480));
    Span4Mux_v I__9932 (
            .O(N__43516),
            .I(N__43477));
    LocalMux I__9931 (
            .O(N__43499),
            .I(N__43470));
    Span4Mux_v I__9930 (
            .O(N__43494),
            .I(N__43470));
    Span4Mux_v I__9929 (
            .O(N__43485),
            .I(N__43470));
    LocalMux I__9928 (
            .O(N__43480),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9927 (
            .O(N__43477),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9926 (
            .O(N__43470),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__9925 (
            .O(N__43463),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3_cascade_ ));
    CascadeMux I__9924 (
            .O(N__43460),
            .I(N__43457));
    InMux I__9923 (
            .O(N__43457),
            .I(N__43453));
    InMux I__9922 (
            .O(N__43456),
            .I(N__43450));
    LocalMux I__9921 (
            .O(N__43453),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    LocalMux I__9920 (
            .O(N__43450),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    InMux I__9919 (
            .O(N__43445),
            .I(N__43442));
    LocalMux I__9918 (
            .O(N__43442),
            .I(N__43431));
    InMux I__9917 (
            .O(N__43441),
            .I(N__43424));
    InMux I__9916 (
            .O(N__43440),
            .I(N__43424));
    InMux I__9915 (
            .O(N__43439),
            .I(N__43424));
    InMux I__9914 (
            .O(N__43438),
            .I(N__43413));
    InMux I__9913 (
            .O(N__43437),
            .I(N__43413));
    InMux I__9912 (
            .O(N__43436),
            .I(N__43413));
    InMux I__9911 (
            .O(N__43435),
            .I(N__43413));
    InMux I__9910 (
            .O(N__43434),
            .I(N__43413));
    Span4Mux_h I__9909 (
            .O(N__43431),
            .I(N__43403));
    LocalMux I__9908 (
            .O(N__43424),
            .I(N__43400));
    LocalMux I__9907 (
            .O(N__43413),
            .I(N__43397));
    InMux I__9906 (
            .O(N__43412),
            .I(N__43382));
    InMux I__9905 (
            .O(N__43411),
            .I(N__43382));
    InMux I__9904 (
            .O(N__43410),
            .I(N__43382));
    InMux I__9903 (
            .O(N__43409),
            .I(N__43382));
    InMux I__9902 (
            .O(N__43408),
            .I(N__43382));
    InMux I__9901 (
            .O(N__43407),
            .I(N__43382));
    InMux I__9900 (
            .O(N__43406),
            .I(N__43382));
    Odrv4 I__9899 (
            .O(N__43403),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    Odrv4 I__9898 (
            .O(N__43400),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    Odrv4 I__9897 (
            .O(N__43397),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    LocalMux I__9896 (
            .O(N__43382),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    CascadeMux I__9895 (
            .O(N__43373),
            .I(N__43370));
    InMux I__9894 (
            .O(N__43370),
            .I(N__43367));
    LocalMux I__9893 (
            .O(N__43367),
            .I(N__43364));
    Span4Mux_h I__9892 (
            .O(N__43364),
            .I(N__43361));
    Odrv4 I__9891 (
            .O(N__43361),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    CEMux I__9890 (
            .O(N__43358),
            .I(N__43355));
    LocalMux I__9889 (
            .O(N__43355),
            .I(N__43349));
    CEMux I__9888 (
            .O(N__43354),
            .I(N__43345));
    CEMux I__9887 (
            .O(N__43353),
            .I(N__43342));
    CEMux I__9886 (
            .O(N__43352),
            .I(N__43339));
    Span4Mux_h I__9885 (
            .O(N__43349),
            .I(N__43336));
    CEMux I__9884 (
            .O(N__43348),
            .I(N__43333));
    LocalMux I__9883 (
            .O(N__43345),
            .I(N__43330));
    LocalMux I__9882 (
            .O(N__43342),
            .I(N__43325));
    LocalMux I__9881 (
            .O(N__43339),
            .I(N__43325));
    Span4Mux_v I__9880 (
            .O(N__43336),
            .I(N__43318));
    LocalMux I__9879 (
            .O(N__43333),
            .I(N__43318));
    Span4Mux_h I__9878 (
            .O(N__43330),
            .I(N__43318));
    Span4Mux_v I__9877 (
            .O(N__43325),
            .I(N__43315));
    Odrv4 I__9876 (
            .O(N__43318),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__9875 (
            .O(N__43315),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__9874 (
            .O(N__43310),
            .I(N__43304));
    InMux I__9873 (
            .O(N__43309),
            .I(N__43304));
    LocalMux I__9872 (
            .O(N__43304),
            .I(N__43293));
    InMux I__9871 (
            .O(N__43303),
            .I(N__43290));
    InMux I__9870 (
            .O(N__43302),
            .I(N__43281));
    InMux I__9869 (
            .O(N__43301),
            .I(N__43281));
    InMux I__9868 (
            .O(N__43300),
            .I(N__43281));
    InMux I__9867 (
            .O(N__43299),
            .I(N__43281));
    InMux I__9866 (
            .O(N__43298),
            .I(N__43274));
    InMux I__9865 (
            .O(N__43297),
            .I(N__43274));
    InMux I__9864 (
            .O(N__43296),
            .I(N__43274));
    Odrv4 I__9863 (
            .O(N__43293),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__9862 (
            .O(N__43290),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__9861 (
            .O(N__43281),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__9860 (
            .O(N__43274),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    InMux I__9859 (
            .O(N__43265),
            .I(N__43260));
    InMux I__9858 (
            .O(N__43264),
            .I(N__43257));
    InMux I__9857 (
            .O(N__43263),
            .I(N__43254));
    LocalMux I__9856 (
            .O(N__43260),
            .I(N__43249));
    LocalMux I__9855 (
            .O(N__43257),
            .I(N__43249));
    LocalMux I__9854 (
            .O(N__43254),
            .I(\phase_controller_inst1.stoper_tr.N_279 ));
    Odrv4 I__9853 (
            .O(N__43249),
            .I(\phase_controller_inst1.stoper_tr.N_279 ));
    InMux I__9852 (
            .O(N__43244),
            .I(N__43238));
    InMux I__9851 (
            .O(N__43243),
            .I(N__43238));
    LocalMux I__9850 (
            .O(N__43238),
            .I(N__43233));
    InMux I__9849 (
            .O(N__43237),
            .I(N__43228));
    InMux I__9848 (
            .O(N__43236),
            .I(N__43228));
    Odrv4 I__9847 (
            .O(N__43233),
            .I(\phase_controller_inst1.stoper_tr.N_262 ));
    LocalMux I__9846 (
            .O(N__43228),
            .I(\phase_controller_inst1.stoper_tr.N_262 ));
    CascadeMux I__9845 (
            .O(N__43223),
            .I(N__43219));
    InMux I__9844 (
            .O(N__43222),
            .I(N__43215));
    InMux I__9843 (
            .O(N__43219),
            .I(N__43212));
    InMux I__9842 (
            .O(N__43218),
            .I(N__43209));
    LocalMux I__9841 (
            .O(N__43215),
            .I(N__43206));
    LocalMux I__9840 (
            .O(N__43212),
            .I(N__43203));
    LocalMux I__9839 (
            .O(N__43209),
            .I(N__43200));
    Span4Mux_v I__9838 (
            .O(N__43206),
            .I(N__43197));
    Odrv12 I__9837 (
            .O(N__43203),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    Odrv4 I__9836 (
            .O(N__43200),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    Odrv4 I__9835 (
            .O(N__43197),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    InMux I__9834 (
            .O(N__43190),
            .I(N__43176));
    InMux I__9833 (
            .O(N__43189),
            .I(N__43176));
    InMux I__9832 (
            .O(N__43188),
            .I(N__43176));
    InMux I__9831 (
            .O(N__43187),
            .I(N__43176));
    InMux I__9830 (
            .O(N__43186),
            .I(N__43171));
    InMux I__9829 (
            .O(N__43185),
            .I(N__43171));
    LocalMux I__9828 (
            .O(N__43176),
            .I(N__43166));
    LocalMux I__9827 (
            .O(N__43171),
            .I(N__43166));
    Span4Mux_h I__9826 (
            .O(N__43166),
            .I(N__43157));
    InMux I__9825 (
            .O(N__43165),
            .I(N__43154));
    InMux I__9824 (
            .O(N__43164),
            .I(N__43143));
    InMux I__9823 (
            .O(N__43163),
            .I(N__43143));
    InMux I__9822 (
            .O(N__43162),
            .I(N__43143));
    InMux I__9821 (
            .O(N__43161),
            .I(N__43143));
    InMux I__9820 (
            .O(N__43160),
            .I(N__43143));
    Odrv4 I__9819 (
            .O(N__43157),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__9818 (
            .O(N__43154),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__9817 (
            .O(N__43143),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    InMux I__9816 (
            .O(N__43136),
            .I(N__43133));
    LocalMux I__9815 (
            .O(N__43133),
            .I(N__43130));
    Span4Mux_h I__9814 (
            .O(N__43130),
            .I(N__43127));
    Odrv4 I__9813 (
            .O(N__43127),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CEMux I__9812 (
            .O(N__43124),
            .I(N__43120));
    CEMux I__9811 (
            .O(N__43123),
            .I(N__43117));
    LocalMux I__9810 (
            .O(N__43120),
            .I(N__43112));
    LocalMux I__9809 (
            .O(N__43117),
            .I(N__43112));
    Span4Mux_v I__9808 (
            .O(N__43112),
            .I(N__43107));
    CEMux I__9807 (
            .O(N__43111),
            .I(N__43104));
    CEMux I__9806 (
            .O(N__43110),
            .I(N__43100));
    Span4Mux_h I__9805 (
            .O(N__43107),
            .I(N__43095));
    LocalMux I__9804 (
            .O(N__43104),
            .I(N__43095));
    CEMux I__9803 (
            .O(N__43103),
            .I(N__43091));
    LocalMux I__9802 (
            .O(N__43100),
            .I(N__43088));
    Span4Mux_v I__9801 (
            .O(N__43095),
            .I(N__43085));
    CEMux I__9800 (
            .O(N__43094),
            .I(N__43082));
    LocalMux I__9799 (
            .O(N__43091),
            .I(N__43079));
    Span4Mux_h I__9798 (
            .O(N__43088),
            .I(N__43076));
    Sp12to4 I__9797 (
            .O(N__43085),
            .I(N__43071));
    LocalMux I__9796 (
            .O(N__43082),
            .I(N__43071));
    Odrv4 I__9795 (
            .O(N__43079),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__9794 (
            .O(N__43076),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__9793 (
            .O(N__43071),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__9792 (
            .O(N__43064),
            .I(N__43058));
    InMux I__9791 (
            .O(N__43063),
            .I(N__43055));
    InMux I__9790 (
            .O(N__43062),
            .I(N__43050));
    InMux I__9789 (
            .O(N__43061),
            .I(N__43050));
    LocalMux I__9788 (
            .O(N__43058),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    LocalMux I__9787 (
            .O(N__43055),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    LocalMux I__9786 (
            .O(N__43050),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    CascadeMux I__9785 (
            .O(N__43043),
            .I(N__43040));
    InMux I__9784 (
            .O(N__43040),
            .I(N__43037));
    LocalMux I__9783 (
            .O(N__43037),
            .I(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__9782 (
            .O(N__43034),
            .I(N__43029));
    InMux I__9781 (
            .O(N__43033),
            .I(N__43024));
    InMux I__9780 (
            .O(N__43032),
            .I(N__43024));
    LocalMux I__9779 (
            .O(N__43029),
            .I(N__43019));
    LocalMux I__9778 (
            .O(N__43024),
            .I(N__43016));
    InMux I__9777 (
            .O(N__43023),
            .I(N__43010));
    InMux I__9776 (
            .O(N__43022),
            .I(N__43010));
    Span4Mux_v I__9775 (
            .O(N__43019),
            .I(N__43007));
    Span4Mux_h I__9774 (
            .O(N__43016),
            .I(N__43004));
    InMux I__9773 (
            .O(N__43015),
            .I(N__43001));
    LocalMux I__9772 (
            .O(N__43010),
            .I(N__42998));
    Odrv4 I__9771 (
            .O(N__43007),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9770 (
            .O(N__43004),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9769 (
            .O(N__43001),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9768 (
            .O(N__42998),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__9767 (
            .O(N__42989),
            .I(N__42985));
    InMux I__9766 (
            .O(N__42988),
            .I(N__42982));
    LocalMux I__9765 (
            .O(N__42985),
            .I(N__42977));
    LocalMux I__9764 (
            .O(N__42982),
            .I(N__42974));
    InMux I__9763 (
            .O(N__42981),
            .I(N__42971));
    InMux I__9762 (
            .O(N__42980),
            .I(N__42968));
    Span12Mux_h I__9761 (
            .O(N__42977),
            .I(N__42965));
    Odrv12 I__9760 (
            .O(N__42974),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__9759 (
            .O(N__42971),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__9758 (
            .O(N__42968),
            .I(\phase_controller_slave.hc_time_passed ));
    Odrv12 I__9757 (
            .O(N__42965),
            .I(\phase_controller_slave.hc_time_passed ));
    InMux I__9756 (
            .O(N__42956),
            .I(N__42953));
    LocalMux I__9755 (
            .O(N__42953),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ));
    CascadeMux I__9754 (
            .O(N__42950),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19_cascade_ ));
    InMux I__9753 (
            .O(N__42947),
            .I(N__42944));
    LocalMux I__9752 (
            .O(N__42944),
            .I(\delay_measurement_inst.delay_tr_timer.N_293 ));
    CascadeMux I__9751 (
            .O(N__42941),
            .I(\delay_measurement_inst.N_358_cascade_ ));
    InMux I__9750 (
            .O(N__42938),
            .I(N__42935));
    LocalMux I__9749 (
            .O(N__42935),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ));
    InMux I__9748 (
            .O(N__42932),
            .I(N__42929));
    LocalMux I__9747 (
            .O(N__42929),
            .I(N__42926));
    Odrv4 I__9746 (
            .O(N__42926),
            .I(\delay_measurement_inst.N_307 ));
    InMux I__9745 (
            .O(N__42923),
            .I(N__42920));
    LocalMux I__9744 (
            .O(N__42920),
            .I(N__42917));
    Span12Mux_h I__9743 (
            .O(N__42917),
            .I(N__42914));
    Odrv12 I__9742 (
            .O(N__42914),
            .I(\phase_controller_slave.start_timer_hc_RNO_0_0 ));
    CascadeMux I__9741 (
            .O(N__42911),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__9740 (
            .O(N__42908),
            .I(N__42905));
    LocalMux I__9739 (
            .O(N__42905),
            .I(N__42900));
    InMux I__9738 (
            .O(N__42904),
            .I(N__42897));
    InMux I__9737 (
            .O(N__42903),
            .I(N__42894));
    Span4Mux_v I__9736 (
            .O(N__42900),
            .I(N__42888));
    LocalMux I__9735 (
            .O(N__42897),
            .I(N__42885));
    LocalMux I__9734 (
            .O(N__42894),
            .I(N__42882));
    InMux I__9733 (
            .O(N__42893),
            .I(N__42877));
    InMux I__9732 (
            .O(N__42892),
            .I(N__42877));
    InMux I__9731 (
            .O(N__42891),
            .I(N__42874));
    Odrv4 I__9730 (
            .O(N__42888),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__9729 (
            .O(N__42885),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__9728 (
            .O(N__42882),
            .I(phase_controller_inst1_state_4));
    LocalMux I__9727 (
            .O(N__42877),
            .I(phase_controller_inst1_state_4));
    LocalMux I__9726 (
            .O(N__42874),
            .I(phase_controller_inst1_state_4));
    InMux I__9725 (
            .O(N__42863),
            .I(N__42856));
    InMux I__9724 (
            .O(N__42862),
            .I(N__42856));
    InMux I__9723 (
            .O(N__42861),
            .I(N__42853));
    LocalMux I__9722 (
            .O(N__42856),
            .I(N__42850));
    LocalMux I__9721 (
            .O(N__42853),
            .I(N__42847));
    Span4Mux_v I__9720 (
            .O(N__42850),
            .I(N__42844));
    Span4Mux_v I__9719 (
            .O(N__42847),
            .I(N__42841));
    Span4Mux_v I__9718 (
            .O(N__42844),
            .I(N__42838));
    Span4Mux_v I__9717 (
            .O(N__42841),
            .I(N__42835));
    Span4Mux_v I__9716 (
            .O(N__42838),
            .I(N__42832));
    Odrv4 I__9715 (
            .O(N__42835),
            .I(il_max_comp2_D2));
    Odrv4 I__9714 (
            .O(N__42832),
            .I(il_max_comp2_D2));
    CascadeMux I__9713 (
            .O(N__42827),
            .I(N__42824));
    InMux I__9712 (
            .O(N__42824),
            .I(N__42818));
    InMux I__9711 (
            .O(N__42823),
            .I(N__42818));
    LocalMux I__9710 (
            .O(N__42818),
            .I(N__42814));
    InMux I__9709 (
            .O(N__42817),
            .I(N__42809));
    Span4Mux_h I__9708 (
            .O(N__42814),
            .I(N__42806));
    InMux I__9707 (
            .O(N__42813),
            .I(N__42803));
    InMux I__9706 (
            .O(N__42812),
            .I(N__42800));
    LocalMux I__9705 (
            .O(N__42809),
            .I(N__42797));
    Span4Mux_h I__9704 (
            .O(N__42806),
            .I(N__42794));
    LocalMux I__9703 (
            .O(N__42803),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__9702 (
            .O(N__42800),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    Odrv4 I__9701 (
            .O(N__42797),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    Odrv4 I__9700 (
            .O(N__42794),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    InMux I__9699 (
            .O(N__42785),
            .I(N__42782));
    LocalMux I__9698 (
            .O(N__42782),
            .I(N__42778));
    InMux I__9697 (
            .O(N__42781),
            .I(N__42775));
    Span4Mux_h I__9696 (
            .O(N__42778),
            .I(N__42771));
    LocalMux I__9695 (
            .O(N__42775),
            .I(N__42768));
    InMux I__9694 (
            .O(N__42774),
            .I(N__42765));
    Span4Mux_v I__9693 (
            .O(N__42771),
            .I(N__42762));
    Odrv12 I__9692 (
            .O(N__42768),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__9691 (
            .O(N__42765),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    Odrv4 I__9690 (
            .O(N__42762),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    InMux I__9689 (
            .O(N__42755),
            .I(bfn_17_16_0_));
    InMux I__9688 (
            .O(N__42752),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__9687 (
            .O(N__42749),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__9686 (
            .O(N__42746),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9685 (
            .O(N__42743),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__9684 (
            .O(N__42740),
            .I(N__42724));
    InMux I__9683 (
            .O(N__42739),
            .I(N__42724));
    InMux I__9682 (
            .O(N__42738),
            .I(N__42724));
    InMux I__9681 (
            .O(N__42737),
            .I(N__42724));
    InMux I__9680 (
            .O(N__42736),
            .I(N__42693));
    InMux I__9679 (
            .O(N__42735),
            .I(N__42693));
    InMux I__9678 (
            .O(N__42734),
            .I(N__42693));
    InMux I__9677 (
            .O(N__42733),
            .I(N__42693));
    LocalMux I__9676 (
            .O(N__42724),
            .I(N__42690));
    InMux I__9675 (
            .O(N__42723),
            .I(N__42681));
    InMux I__9674 (
            .O(N__42722),
            .I(N__42681));
    InMux I__9673 (
            .O(N__42721),
            .I(N__42681));
    InMux I__9672 (
            .O(N__42720),
            .I(N__42681));
    InMux I__9671 (
            .O(N__42719),
            .I(N__42672));
    InMux I__9670 (
            .O(N__42718),
            .I(N__42672));
    InMux I__9669 (
            .O(N__42717),
            .I(N__42672));
    InMux I__9668 (
            .O(N__42716),
            .I(N__42672));
    InMux I__9667 (
            .O(N__42715),
            .I(N__42663));
    InMux I__9666 (
            .O(N__42714),
            .I(N__42663));
    InMux I__9665 (
            .O(N__42713),
            .I(N__42663));
    InMux I__9664 (
            .O(N__42712),
            .I(N__42663));
    InMux I__9663 (
            .O(N__42711),
            .I(N__42654));
    InMux I__9662 (
            .O(N__42710),
            .I(N__42654));
    InMux I__9661 (
            .O(N__42709),
            .I(N__42654));
    InMux I__9660 (
            .O(N__42708),
            .I(N__42654));
    InMux I__9659 (
            .O(N__42707),
            .I(N__42649));
    InMux I__9658 (
            .O(N__42706),
            .I(N__42649));
    InMux I__9657 (
            .O(N__42705),
            .I(N__42640));
    InMux I__9656 (
            .O(N__42704),
            .I(N__42640));
    InMux I__9655 (
            .O(N__42703),
            .I(N__42640));
    InMux I__9654 (
            .O(N__42702),
            .I(N__42640));
    LocalMux I__9653 (
            .O(N__42693),
            .I(N__42633));
    Span4Mux_h I__9652 (
            .O(N__42690),
            .I(N__42633));
    LocalMux I__9651 (
            .O(N__42681),
            .I(N__42633));
    LocalMux I__9650 (
            .O(N__42672),
            .I(N__42626));
    LocalMux I__9649 (
            .O(N__42663),
            .I(N__42626));
    LocalMux I__9648 (
            .O(N__42654),
            .I(N__42626));
    LocalMux I__9647 (
            .O(N__42649),
            .I(N__42621));
    LocalMux I__9646 (
            .O(N__42640),
            .I(N__42621));
    Span4Mux_v I__9645 (
            .O(N__42633),
            .I(N__42616));
    Span4Mux_v I__9644 (
            .O(N__42626),
            .I(N__42616));
    Span4Mux_h I__9643 (
            .O(N__42621),
            .I(N__42613));
    Span4Mux_h I__9642 (
            .O(N__42616),
            .I(N__42610));
    Span4Mux_v I__9641 (
            .O(N__42613),
            .I(N__42607));
    Odrv4 I__9640 (
            .O(N__42610),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9639 (
            .O(N__42607),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9638 (
            .O(N__42602),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__9637 (
            .O(N__42599),
            .I(N__42596));
    LocalMux I__9636 (
            .O(N__42596),
            .I(N__42592));
    CEMux I__9635 (
            .O(N__42595),
            .I(N__42587));
    Span4Mux_h I__9634 (
            .O(N__42592),
            .I(N__42584));
    CEMux I__9633 (
            .O(N__42591),
            .I(N__42581));
    CEMux I__9632 (
            .O(N__42590),
            .I(N__42578));
    LocalMux I__9631 (
            .O(N__42587),
            .I(N__42575));
    Span4Mux_h I__9630 (
            .O(N__42584),
            .I(N__42572));
    LocalMux I__9629 (
            .O(N__42581),
            .I(N__42569));
    LocalMux I__9628 (
            .O(N__42578),
            .I(N__42566));
    Span4Mux_v I__9627 (
            .O(N__42575),
            .I(N__42563));
    Sp12to4 I__9626 (
            .O(N__42572),
            .I(N__42560));
    Span4Mux_h I__9625 (
            .O(N__42569),
            .I(N__42557));
    Span4Mux_h I__9624 (
            .O(N__42566),
            .I(N__42554));
    Span4Mux_v I__9623 (
            .O(N__42563),
            .I(N__42551));
    Span12Mux_v I__9622 (
            .O(N__42560),
            .I(N__42548));
    Span4Mux_v I__9621 (
            .O(N__42557),
            .I(N__42545));
    Span4Mux_v I__9620 (
            .O(N__42554),
            .I(N__42542));
    Odrv4 I__9619 (
            .O(N__42551),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv12 I__9618 (
            .O(N__42548),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv4 I__9617 (
            .O(N__42545),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv4 I__9616 (
            .O(N__42542),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    InMux I__9615 (
            .O(N__42533),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__9614 (
            .O(N__42530),
            .I(bfn_17_15_0_));
    InMux I__9613 (
            .O(N__42527),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__9612 (
            .O(N__42524),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__9611 (
            .O(N__42521),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__9610 (
            .O(N__42518),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__9609 (
            .O(N__42515),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__9608 (
            .O(N__42512),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__9607 (
            .O(N__42509),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9606 (
            .O(N__42506),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__9605 (
            .O(N__42503),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__9604 (
            .O(N__42500),
            .I(bfn_17_14_0_));
    InMux I__9603 (
            .O(N__42497),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__9602 (
            .O(N__42494),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__9601 (
            .O(N__42491),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__9600 (
            .O(N__42488),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__9599 (
            .O(N__42485),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__9598 (
            .O(N__42482),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__9597 (
            .O(N__42479),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__9596 (
            .O(N__42476),
            .I(N__42471));
    InMux I__9595 (
            .O(N__42475),
            .I(N__42467));
    InMux I__9594 (
            .O(N__42474),
            .I(N__42464));
    LocalMux I__9593 (
            .O(N__42471),
            .I(N__42461));
    InMux I__9592 (
            .O(N__42470),
            .I(N__42458));
    LocalMux I__9591 (
            .O(N__42467),
            .I(N__42455));
    LocalMux I__9590 (
            .O(N__42464),
            .I(N__42448));
    Span4Mux_h I__9589 (
            .O(N__42461),
            .I(N__42448));
    LocalMux I__9588 (
            .O(N__42458),
            .I(N__42448));
    Span4Mux_h I__9587 (
            .O(N__42455),
            .I(N__42445));
    Span4Mux_v I__9586 (
            .O(N__42448),
            .I(N__42442));
    Odrv4 I__9585 (
            .O(N__42445),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    Odrv4 I__9584 (
            .O(N__42442),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__9583 (
            .O(N__42437),
            .I(N__42433));
    InMux I__9582 (
            .O(N__42436),
            .I(N__42428));
    LocalMux I__9581 (
            .O(N__42433),
            .I(N__42425));
    InMux I__9580 (
            .O(N__42432),
            .I(N__42422));
    InMux I__9579 (
            .O(N__42431),
            .I(N__42419));
    LocalMux I__9578 (
            .O(N__42428),
            .I(N__42416));
    Span4Mux_h I__9577 (
            .O(N__42425),
            .I(N__42409));
    LocalMux I__9576 (
            .O(N__42422),
            .I(N__42409));
    LocalMux I__9575 (
            .O(N__42419),
            .I(N__42409));
    Span4Mux_h I__9574 (
            .O(N__42416),
            .I(N__42404));
    Span4Mux_v I__9573 (
            .O(N__42409),
            .I(N__42404));
    Odrv4 I__9572 (
            .O(N__42404),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    CascadeMux I__9571 (
            .O(N__42401),
            .I(N__42398));
    InMux I__9570 (
            .O(N__42398),
            .I(N__42395));
    LocalMux I__9569 (
            .O(N__42395),
            .I(N__42392));
    Span4Mux_h I__9568 (
            .O(N__42392),
            .I(N__42388));
    InMux I__9567 (
            .O(N__42391),
            .I(N__42385));
    Odrv4 I__9566 (
            .O(N__42388),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2 ));
    LocalMux I__9565 (
            .O(N__42385),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2 ));
    CascadeMux I__9564 (
            .O(N__42380),
            .I(N__42376));
    InMux I__9563 (
            .O(N__42379),
            .I(N__42373));
    InMux I__9562 (
            .O(N__42376),
            .I(N__42370));
    LocalMux I__9561 (
            .O(N__42373),
            .I(N__42366));
    LocalMux I__9560 (
            .O(N__42370),
            .I(N__42363));
    InMux I__9559 (
            .O(N__42369),
            .I(N__42360));
    Span4Mux_h I__9558 (
            .O(N__42366),
            .I(N__42357));
    Span12Mux_v I__9557 (
            .O(N__42363),
            .I(N__42354));
    LocalMux I__9556 (
            .O(N__42360),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    Odrv4 I__9555 (
            .O(N__42357),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    Odrv12 I__9554 (
            .O(N__42354),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    CascadeMux I__9553 (
            .O(N__42347),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4Z0Z_3_cascade_ ));
    InMux I__9552 (
            .O(N__42344),
            .I(N__42341));
    LocalMux I__9551 (
            .O(N__42341),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_7_0 ));
    InMux I__9550 (
            .O(N__42338),
            .I(bfn_17_13_0_));
    InMux I__9549 (
            .O(N__42335),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__9548 (
            .O(N__42332),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__9547 (
            .O(N__42329),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__9546 (
            .O(N__42326),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__9545 (
            .O(N__42323),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__9544 (
            .O(N__42320),
            .I(N__42315));
    InMux I__9543 (
            .O(N__42319),
            .I(N__42312));
    InMux I__9542 (
            .O(N__42318),
            .I(N__42309));
    InMux I__9541 (
            .O(N__42315),
            .I(N__42306));
    LocalMux I__9540 (
            .O(N__42312),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__9539 (
            .O(N__42309),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__9538 (
            .O(N__42306),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__9537 (
            .O(N__42299),
            .I(N__42296));
    LocalMux I__9536 (
            .O(N__42296),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__9535 (
            .O(N__42293),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__9534 (
            .O(N__42290),
            .I(N__42285));
    InMux I__9533 (
            .O(N__42289),
            .I(N__42282));
    InMux I__9532 (
            .O(N__42288),
            .I(N__42279));
    InMux I__9531 (
            .O(N__42285),
            .I(N__42276));
    LocalMux I__9530 (
            .O(N__42282),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__9529 (
            .O(N__42279),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__9528 (
            .O(N__42276),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__9527 (
            .O(N__42269),
            .I(N__42266));
    LocalMux I__9526 (
            .O(N__42266),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__9525 (
            .O(N__42263),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__9524 (
            .O(N__42260),
            .I(N__42255));
    InMux I__9523 (
            .O(N__42259),
            .I(N__42252));
    InMux I__9522 (
            .O(N__42258),
            .I(N__42249));
    InMux I__9521 (
            .O(N__42255),
            .I(N__42246));
    LocalMux I__9520 (
            .O(N__42252),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__9519 (
            .O(N__42249),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__9518 (
            .O(N__42246),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__9517 (
            .O(N__42239),
            .I(N__42236));
    LocalMux I__9516 (
            .O(N__42236),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__9515 (
            .O(N__42233),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__9514 (
            .O(N__42230),
            .I(N__42225));
    InMux I__9513 (
            .O(N__42229),
            .I(N__42222));
    InMux I__9512 (
            .O(N__42228),
            .I(N__42219));
    InMux I__9511 (
            .O(N__42225),
            .I(N__42216));
    LocalMux I__9510 (
            .O(N__42222),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__9509 (
            .O(N__42219),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__9508 (
            .O(N__42216),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__9507 (
            .O(N__42209),
            .I(N__42206));
    LocalMux I__9506 (
            .O(N__42206),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__9505 (
            .O(N__42203),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__9504 (
            .O(N__42200),
            .I(N__42195));
    InMux I__9503 (
            .O(N__42199),
            .I(N__42192));
    InMux I__9502 (
            .O(N__42198),
            .I(N__42189));
    InMux I__9501 (
            .O(N__42195),
            .I(N__42186));
    LocalMux I__9500 (
            .O(N__42192),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__9499 (
            .O(N__42189),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__9498 (
            .O(N__42186),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__9497 (
            .O(N__42179),
            .I(N__42176));
    LocalMux I__9496 (
            .O(N__42176),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__9495 (
            .O(N__42173),
            .I(bfn_17_11_0_));
    CascadeMux I__9494 (
            .O(N__42170),
            .I(N__42165));
    InMux I__9493 (
            .O(N__42169),
            .I(N__42162));
    InMux I__9492 (
            .O(N__42168),
            .I(N__42159));
    InMux I__9491 (
            .O(N__42165),
            .I(N__42156));
    LocalMux I__9490 (
            .O(N__42162),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__9489 (
            .O(N__42159),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__9488 (
            .O(N__42156),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__9487 (
            .O(N__42149),
            .I(N__42146));
    LocalMux I__9486 (
            .O(N__42146),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__9485 (
            .O(N__42143),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__9484 (
            .O(N__42140),
            .I(N__42135));
    InMux I__9483 (
            .O(N__42139),
            .I(N__42132));
    InMux I__9482 (
            .O(N__42138),
            .I(N__42129));
    InMux I__9481 (
            .O(N__42135),
            .I(N__42126));
    LocalMux I__9480 (
            .O(N__42132),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__9479 (
            .O(N__42129),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__9478 (
            .O(N__42126),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    CascadeMux I__9477 (
            .O(N__42119),
            .I(N__42115));
    InMux I__9476 (
            .O(N__42118),
            .I(N__42112));
    InMux I__9475 (
            .O(N__42115),
            .I(N__42109));
    LocalMux I__9474 (
            .O(N__42112),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__9473 (
            .O(N__42109),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__9472 (
            .O(N__42104),
            .I(N__42101));
    LocalMux I__9471 (
            .O(N__42101),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__9470 (
            .O(N__42098),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__9469 (
            .O(N__42095),
            .I(N__42090));
    InMux I__9468 (
            .O(N__42094),
            .I(N__42087));
    InMux I__9467 (
            .O(N__42093),
            .I(N__42084));
    InMux I__9466 (
            .O(N__42090),
            .I(N__42081));
    LocalMux I__9465 (
            .O(N__42087),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__9464 (
            .O(N__42084),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__9463 (
            .O(N__42081),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    CascadeMux I__9462 (
            .O(N__42074),
            .I(N__42070));
    InMux I__9461 (
            .O(N__42073),
            .I(N__42067));
    InMux I__9460 (
            .O(N__42070),
            .I(N__42064));
    LocalMux I__9459 (
            .O(N__42067),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__9458 (
            .O(N__42064),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__9457 (
            .O(N__42059),
            .I(N__42056));
    InMux I__9456 (
            .O(N__42056),
            .I(N__42053));
    LocalMux I__9455 (
            .O(N__42053),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ));
    InMux I__9454 (
            .O(N__42050),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    CascadeMux I__9453 (
            .O(N__42047),
            .I(N__42042));
    InMux I__9452 (
            .O(N__42046),
            .I(N__42039));
    InMux I__9451 (
            .O(N__42045),
            .I(N__42036));
    InMux I__9450 (
            .O(N__42042),
            .I(N__42033));
    LocalMux I__9449 (
            .O(N__42039),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__9448 (
            .O(N__42036),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__9447 (
            .O(N__42033),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__9446 (
            .O(N__42026),
            .I(N__42023));
    LocalMux I__9445 (
            .O(N__42023),
            .I(N__42020));
    Span4Mux_h I__9444 (
            .O(N__42020),
            .I(N__42017));
    Span4Mux_h I__9443 (
            .O(N__42017),
            .I(N__42013));
    CascadeMux I__9442 (
            .O(N__42016),
            .I(N__42007));
    Span4Mux_v I__9441 (
            .O(N__42013),
            .I(N__42004));
    InMux I__9440 (
            .O(N__42012),
            .I(N__42001));
    InMux I__9439 (
            .O(N__42011),
            .I(N__41998));
    CascadeMux I__9438 (
            .O(N__42010),
            .I(N__41995));
    InMux I__9437 (
            .O(N__42007),
            .I(N__41992));
    Span4Mux_h I__9436 (
            .O(N__42004),
            .I(N__41987));
    LocalMux I__9435 (
            .O(N__42001),
            .I(N__41987));
    LocalMux I__9434 (
            .O(N__41998),
            .I(N__41984));
    InMux I__9433 (
            .O(N__41995),
            .I(N__41981));
    LocalMux I__9432 (
            .O(N__41992),
            .I(N__41978));
    Span4Mux_v I__9431 (
            .O(N__41987),
            .I(N__41975));
    Span4Mux_v I__9430 (
            .O(N__41984),
            .I(N__41970));
    LocalMux I__9429 (
            .O(N__41981),
            .I(N__41970));
    Odrv12 I__9428 (
            .O(N__41978),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__9427 (
            .O(N__41975),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__9426 (
            .O(N__41970),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__9425 (
            .O(N__41963),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__9424 (
            .O(N__41960),
            .I(N__41955));
    InMux I__9423 (
            .O(N__41959),
            .I(N__41952));
    InMux I__9422 (
            .O(N__41958),
            .I(N__41949));
    InMux I__9421 (
            .O(N__41955),
            .I(N__41946));
    LocalMux I__9420 (
            .O(N__41952),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__9419 (
            .O(N__41949),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__9418 (
            .O(N__41946),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__9417 (
            .O(N__41939),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__9416 (
            .O(N__41936),
            .I(N__41931));
    InMux I__9415 (
            .O(N__41935),
            .I(N__41928));
    InMux I__9414 (
            .O(N__41934),
            .I(N__41925));
    InMux I__9413 (
            .O(N__41931),
            .I(N__41922));
    LocalMux I__9412 (
            .O(N__41928),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__9411 (
            .O(N__41925),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__9410 (
            .O(N__41922),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__9409 (
            .O(N__41915),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__9408 (
            .O(N__41912),
            .I(N__41907));
    InMux I__9407 (
            .O(N__41911),
            .I(N__41904));
    InMux I__9406 (
            .O(N__41910),
            .I(N__41901));
    InMux I__9405 (
            .O(N__41907),
            .I(N__41898));
    LocalMux I__9404 (
            .O(N__41904),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__9403 (
            .O(N__41901),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__9402 (
            .O(N__41898),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__9401 (
            .O(N__41891),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__9400 (
            .O(N__41888),
            .I(N__41883));
    InMux I__9399 (
            .O(N__41887),
            .I(N__41880));
    InMux I__9398 (
            .O(N__41886),
            .I(N__41877));
    InMux I__9397 (
            .O(N__41883),
            .I(N__41874));
    LocalMux I__9396 (
            .O(N__41880),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__9395 (
            .O(N__41877),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__9394 (
            .O(N__41874),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__9393 (
            .O(N__41867),
            .I(bfn_17_10_0_));
    CascadeMux I__9392 (
            .O(N__41864),
            .I(N__41859));
    InMux I__9391 (
            .O(N__41863),
            .I(N__41856));
    InMux I__9390 (
            .O(N__41862),
            .I(N__41853));
    InMux I__9389 (
            .O(N__41859),
            .I(N__41850));
    LocalMux I__9388 (
            .O(N__41856),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__9387 (
            .O(N__41853),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__9386 (
            .O(N__41850),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    CascadeMux I__9385 (
            .O(N__41843),
            .I(N__41840));
    InMux I__9384 (
            .O(N__41840),
            .I(N__41837));
    LocalMux I__9383 (
            .O(N__41837),
            .I(N__41833));
    InMux I__9382 (
            .O(N__41836),
            .I(N__41830));
    Odrv4 I__9381 (
            .O(N__41833),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__9380 (
            .O(N__41830),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__9379 (
            .O(N__41825),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__9378 (
            .O(N__41822),
            .I(N__41817));
    InMux I__9377 (
            .O(N__41821),
            .I(N__41814));
    InMux I__9376 (
            .O(N__41820),
            .I(N__41811));
    InMux I__9375 (
            .O(N__41817),
            .I(N__41808));
    LocalMux I__9374 (
            .O(N__41814),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__9373 (
            .O(N__41811),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__9372 (
            .O(N__41808),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__9371 (
            .O(N__41801),
            .I(N__41798));
    LocalMux I__9370 (
            .O(N__41798),
            .I(N__41794));
    InMux I__9369 (
            .O(N__41797),
            .I(N__41791));
    Span4Mux_v I__9368 (
            .O(N__41794),
            .I(N__41788));
    LocalMux I__9367 (
            .O(N__41791),
            .I(N__41785));
    Odrv4 I__9366 (
            .O(N__41788),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__9365 (
            .O(N__41785),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__9364 (
            .O(N__41780),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__9363 (
            .O(N__41777),
            .I(N__41772));
    InMux I__9362 (
            .O(N__41776),
            .I(N__41769));
    InMux I__9361 (
            .O(N__41775),
            .I(N__41766));
    InMux I__9360 (
            .O(N__41772),
            .I(N__41763));
    LocalMux I__9359 (
            .O(N__41769),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__9358 (
            .O(N__41766),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__9357 (
            .O(N__41763),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__9356 (
            .O(N__41756),
            .I(N__41753));
    LocalMux I__9355 (
            .O(N__41753),
            .I(N__41749));
    CascadeMux I__9354 (
            .O(N__41752),
            .I(N__41746));
    Span4Mux_v I__9353 (
            .O(N__41749),
            .I(N__41743));
    InMux I__9352 (
            .O(N__41746),
            .I(N__41740));
    Odrv4 I__9351 (
            .O(N__41743),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__9350 (
            .O(N__41740),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__9349 (
            .O(N__41735),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__9348 (
            .O(N__41732),
            .I(N__41727));
    InMux I__9347 (
            .O(N__41731),
            .I(N__41724));
    InMux I__9346 (
            .O(N__41730),
            .I(N__41721));
    InMux I__9345 (
            .O(N__41727),
            .I(N__41718));
    LocalMux I__9344 (
            .O(N__41724),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__9343 (
            .O(N__41721),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__9342 (
            .O(N__41718),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    CascadeMux I__9341 (
            .O(N__41711),
            .I(N__41708));
    InMux I__9340 (
            .O(N__41708),
            .I(N__41702));
    InMux I__9339 (
            .O(N__41707),
            .I(N__41699));
    InMux I__9338 (
            .O(N__41706),
            .I(N__41693));
    InMux I__9337 (
            .O(N__41705),
            .I(N__41693));
    LocalMux I__9336 (
            .O(N__41702),
            .I(N__41688));
    LocalMux I__9335 (
            .O(N__41699),
            .I(N__41688));
    InMux I__9334 (
            .O(N__41698),
            .I(N__41685));
    LocalMux I__9333 (
            .O(N__41693),
            .I(N__41682));
    Span4Mux_v I__9332 (
            .O(N__41688),
            .I(N__41679));
    LocalMux I__9331 (
            .O(N__41685),
            .I(N__41674));
    Span4Mux_h I__9330 (
            .O(N__41682),
            .I(N__41674));
    Odrv4 I__9329 (
            .O(N__41679),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    Odrv4 I__9328 (
            .O(N__41674),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__9327 (
            .O(N__41669),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9326 (
            .O(N__41666),
            .I(N__41661));
    InMux I__9325 (
            .O(N__41665),
            .I(N__41658));
    InMux I__9324 (
            .O(N__41664),
            .I(N__41655));
    InMux I__9323 (
            .O(N__41661),
            .I(N__41652));
    LocalMux I__9322 (
            .O(N__41658),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__9321 (
            .O(N__41655),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__9320 (
            .O(N__41652),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    CascadeMux I__9319 (
            .O(N__41645),
            .I(N__41639));
    InMux I__9318 (
            .O(N__41644),
            .I(N__41635));
    InMux I__9317 (
            .O(N__41643),
            .I(N__41632));
    InMux I__9316 (
            .O(N__41642),
            .I(N__41629));
    InMux I__9315 (
            .O(N__41639),
            .I(N__41624));
    InMux I__9314 (
            .O(N__41638),
            .I(N__41624));
    LocalMux I__9313 (
            .O(N__41635),
            .I(N__41619));
    LocalMux I__9312 (
            .O(N__41632),
            .I(N__41619));
    LocalMux I__9311 (
            .O(N__41629),
            .I(N__41614));
    LocalMux I__9310 (
            .O(N__41624),
            .I(N__41614));
    Span4Mux_v I__9309 (
            .O(N__41619),
            .I(N__41611));
    Span4Mux_h I__9308 (
            .O(N__41614),
            .I(N__41608));
    Odrv4 I__9307 (
            .O(N__41611),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    Odrv4 I__9306 (
            .O(N__41608),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__9305 (
            .O(N__41603),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__9304 (
            .O(N__41600),
            .I(N__41595));
    InMux I__9303 (
            .O(N__41599),
            .I(N__41592));
    InMux I__9302 (
            .O(N__41598),
            .I(N__41589));
    InMux I__9301 (
            .O(N__41595),
            .I(N__41586));
    LocalMux I__9300 (
            .O(N__41592),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__9299 (
            .O(N__41589),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__9298 (
            .O(N__41586),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__9297 (
            .O(N__41579),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__9296 (
            .O(N__41576),
            .I(N__41571));
    InMux I__9295 (
            .O(N__41575),
            .I(N__41568));
    InMux I__9294 (
            .O(N__41574),
            .I(N__41565));
    InMux I__9293 (
            .O(N__41571),
            .I(N__41562));
    LocalMux I__9292 (
            .O(N__41568),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__9291 (
            .O(N__41565),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__9290 (
            .O(N__41562),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    CascadeMux I__9289 (
            .O(N__41555),
            .I(N__41551));
    CascadeMux I__9288 (
            .O(N__41554),
            .I(N__41547));
    InMux I__9287 (
            .O(N__41551),
            .I(N__41544));
    InMux I__9286 (
            .O(N__41550),
            .I(N__41541));
    InMux I__9285 (
            .O(N__41547),
            .I(N__41538));
    LocalMux I__9284 (
            .O(N__41544),
            .I(N__41535));
    LocalMux I__9283 (
            .O(N__41541),
            .I(N__41530));
    LocalMux I__9282 (
            .O(N__41538),
            .I(N__41530));
    Span4Mux_h I__9281 (
            .O(N__41535),
            .I(N__41527));
    Span4Mux_h I__9280 (
            .O(N__41530),
            .I(N__41524));
    Odrv4 I__9279 (
            .O(N__41527),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    Odrv4 I__9278 (
            .O(N__41524),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__9277 (
            .O(N__41519),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__9276 (
            .O(N__41516),
            .I(N__41511));
    InMux I__9275 (
            .O(N__41515),
            .I(N__41508));
    InMux I__9274 (
            .O(N__41514),
            .I(N__41505));
    InMux I__9273 (
            .O(N__41511),
            .I(N__41502));
    LocalMux I__9272 (
            .O(N__41508),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__9271 (
            .O(N__41505),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__9270 (
            .O(N__41502),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    CascadeMux I__9269 (
            .O(N__41495),
            .I(N__41492));
    InMux I__9268 (
            .O(N__41492),
            .I(N__41489));
    LocalMux I__9267 (
            .O(N__41489),
            .I(N__41484));
    InMux I__9266 (
            .O(N__41488),
            .I(N__41479));
    InMux I__9265 (
            .O(N__41487),
            .I(N__41479));
    Span12Mux_v I__9264 (
            .O(N__41484),
            .I(N__41474));
    LocalMux I__9263 (
            .O(N__41479),
            .I(N__41474));
    Odrv12 I__9262 (
            .O(N__41474),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__9261 (
            .O(N__41471),
            .I(bfn_17_9_0_));
    CascadeMux I__9260 (
            .O(N__41468),
            .I(N__41463));
    InMux I__9259 (
            .O(N__41467),
            .I(N__41460));
    InMux I__9258 (
            .O(N__41466),
            .I(N__41457));
    InMux I__9257 (
            .O(N__41463),
            .I(N__41454));
    LocalMux I__9256 (
            .O(N__41460),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__9255 (
            .O(N__41457),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__9254 (
            .O(N__41454),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__9253 (
            .O(N__41447),
            .I(N__41443));
    CascadeMux I__9252 (
            .O(N__41446),
            .I(N__41439));
    LocalMux I__9251 (
            .O(N__41443),
            .I(N__41436));
    InMux I__9250 (
            .O(N__41442),
            .I(N__41431));
    InMux I__9249 (
            .O(N__41439),
            .I(N__41431));
    Span4Mux_v I__9248 (
            .O(N__41436),
            .I(N__41428));
    LocalMux I__9247 (
            .O(N__41431),
            .I(N__41425));
    Odrv4 I__9246 (
            .O(N__41428),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    Odrv12 I__9245 (
            .O(N__41425),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__9244 (
            .O(N__41420),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__9243 (
            .O(N__41417),
            .I(N__41412));
    InMux I__9242 (
            .O(N__41416),
            .I(N__41409));
    InMux I__9241 (
            .O(N__41415),
            .I(N__41406));
    InMux I__9240 (
            .O(N__41412),
            .I(N__41403));
    LocalMux I__9239 (
            .O(N__41409),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__9238 (
            .O(N__41406),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__9237 (
            .O(N__41403),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    CascadeMux I__9236 (
            .O(N__41396),
            .I(N__41392));
    CascadeMux I__9235 (
            .O(N__41395),
            .I(N__41388));
    InMux I__9234 (
            .O(N__41392),
            .I(N__41385));
    InMux I__9233 (
            .O(N__41391),
            .I(N__41380));
    InMux I__9232 (
            .O(N__41388),
            .I(N__41380));
    LocalMux I__9231 (
            .O(N__41385),
            .I(N__41377));
    LocalMux I__9230 (
            .O(N__41380),
            .I(N__41374));
    Span4Mux_h I__9229 (
            .O(N__41377),
            .I(N__41369));
    Span4Mux_h I__9228 (
            .O(N__41374),
            .I(N__41369));
    Odrv4 I__9227 (
            .O(N__41369),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__9226 (
            .O(N__41366),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__9225 (
            .O(N__41363),
            .I(N__41358));
    InMux I__9224 (
            .O(N__41362),
            .I(N__41355));
    InMux I__9223 (
            .O(N__41361),
            .I(N__41352));
    InMux I__9222 (
            .O(N__41358),
            .I(N__41349));
    LocalMux I__9221 (
            .O(N__41355),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__9220 (
            .O(N__41352),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__9219 (
            .O(N__41349),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__9218 (
            .O(N__41342),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__9217 (
            .O(N__41339),
            .I(N__41336));
    InMux I__9216 (
            .O(N__41336),
            .I(N__41333));
    LocalMux I__9215 (
            .O(N__41333),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__9214 (
            .O(N__41330),
            .I(N__41327));
    InMux I__9213 (
            .O(N__41327),
            .I(N__41324));
    LocalMux I__9212 (
            .O(N__41324),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__9211 (
            .O(N__41321),
            .I(N__41318));
    InMux I__9210 (
            .O(N__41318),
            .I(N__41315));
    LocalMux I__9209 (
            .O(N__41315),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__9208 (
            .O(N__41312),
            .I(N__41308));
    InMux I__9207 (
            .O(N__41311),
            .I(N__41305));
    LocalMux I__9206 (
            .O(N__41308),
            .I(N__41301));
    LocalMux I__9205 (
            .O(N__41305),
            .I(N__41298));
    InMux I__9204 (
            .O(N__41304),
            .I(N__41295));
    Odrv12 I__9203 (
            .O(N__41301),
            .I(measured_delay_tr_12));
    Odrv4 I__9202 (
            .O(N__41298),
            .I(measured_delay_tr_12));
    LocalMux I__9201 (
            .O(N__41295),
            .I(measured_delay_tr_12));
    CascadeMux I__9200 (
            .O(N__41288),
            .I(N__41285));
    InMux I__9199 (
            .O(N__41285),
            .I(N__41282));
    LocalMux I__9198 (
            .O(N__41282),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__9197 (
            .O(N__41279),
            .I(N__41276));
    LocalMux I__9196 (
            .O(N__41276),
            .I(N__41273));
    Span4Mux_v I__9195 (
            .O(N__41273),
            .I(N__41269));
    InMux I__9194 (
            .O(N__41272),
            .I(N__41266));
    Span4Mux_h I__9193 (
            .O(N__41269),
            .I(N__41263));
    LocalMux I__9192 (
            .O(N__41266),
            .I(N__41260));
    Span4Mux_h I__9191 (
            .O(N__41263),
            .I(N__41257));
    Span4Mux_v I__9190 (
            .O(N__41260),
            .I(N__41254));
    Odrv4 I__9189 (
            .O(N__41257),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    Odrv4 I__9188 (
            .O(N__41254),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    InMux I__9187 (
            .O(N__41249),
            .I(N__41244));
    InMux I__9186 (
            .O(N__41248),
            .I(N__41241));
    InMux I__9185 (
            .O(N__41247),
            .I(N__41238));
    LocalMux I__9184 (
            .O(N__41244),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9183 (
            .O(N__41241),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9182 (
            .O(N__41238),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__9181 (
            .O(N__41231),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__9180 (
            .O(N__41228),
            .I(N__41223));
    InMux I__9179 (
            .O(N__41227),
            .I(N__41220));
    InMux I__9178 (
            .O(N__41226),
            .I(N__41217));
    InMux I__9177 (
            .O(N__41223),
            .I(N__41214));
    LocalMux I__9176 (
            .O(N__41220),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__9175 (
            .O(N__41217),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__9174 (
            .O(N__41214),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__9173 (
            .O(N__41207),
            .I(N__41202));
    InMux I__9172 (
            .O(N__41206),
            .I(N__41199));
    InMux I__9171 (
            .O(N__41205),
            .I(N__41196));
    LocalMux I__9170 (
            .O(N__41202),
            .I(N__41193));
    LocalMux I__9169 (
            .O(N__41199),
            .I(N__41190));
    LocalMux I__9168 (
            .O(N__41196),
            .I(N__41187));
    Span4Mux_h I__9167 (
            .O(N__41193),
            .I(N__41184));
    Span4Mux_h I__9166 (
            .O(N__41190),
            .I(N__41181));
    Odrv4 I__9165 (
            .O(N__41187),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    Odrv4 I__9164 (
            .O(N__41184),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    Odrv4 I__9163 (
            .O(N__41181),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__9162 (
            .O(N__41174),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__9161 (
            .O(N__41171),
            .I(N__41166));
    InMux I__9160 (
            .O(N__41170),
            .I(N__41163));
    InMux I__9159 (
            .O(N__41169),
            .I(N__41160));
    InMux I__9158 (
            .O(N__41166),
            .I(N__41157));
    LocalMux I__9157 (
            .O(N__41163),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__9156 (
            .O(N__41160),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__9155 (
            .O(N__41157),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__9154 (
            .O(N__41150),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__9153 (
            .O(N__41147),
            .I(N__41144));
    LocalMux I__9152 (
            .O(N__41144),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__9151 (
            .O(N__41141),
            .I(N__41138));
    InMux I__9150 (
            .O(N__41138),
            .I(N__41135));
    LocalMux I__9149 (
            .O(N__41135),
            .I(N__41132));
    Odrv4 I__9148 (
            .O(N__41132),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__9147 (
            .O(N__41129),
            .I(N__41126));
    InMux I__9146 (
            .O(N__41126),
            .I(N__41123));
    LocalMux I__9145 (
            .O(N__41123),
            .I(N__41120));
    Span4Mux_h I__9144 (
            .O(N__41120),
            .I(N__41117));
    Odrv4 I__9143 (
            .O(N__41117),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__9142 (
            .O(N__41114),
            .I(N__41111));
    InMux I__9141 (
            .O(N__41111),
            .I(N__41108));
    LocalMux I__9140 (
            .O(N__41108),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__9139 (
            .O(N__41105),
            .I(N__41102));
    InMux I__9138 (
            .O(N__41102),
            .I(N__41099));
    LocalMux I__9137 (
            .O(N__41099),
            .I(N__41096));
    Span4Mux_v I__9136 (
            .O(N__41096),
            .I(N__41093));
    Odrv4 I__9135 (
            .O(N__41093),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__9134 (
            .O(N__41090),
            .I(N__41087));
    InMux I__9133 (
            .O(N__41087),
            .I(N__41084));
    LocalMux I__9132 (
            .O(N__41084),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__9131 (
            .O(N__41081),
            .I(N__41077));
    InMux I__9130 (
            .O(N__41080),
            .I(N__41074));
    LocalMux I__9129 (
            .O(N__41077),
            .I(N__41070));
    LocalMux I__9128 (
            .O(N__41074),
            .I(N__41067));
    InMux I__9127 (
            .O(N__41073),
            .I(N__41064));
    Odrv12 I__9126 (
            .O(N__41070),
            .I(measured_delay_tr_10));
    Odrv4 I__9125 (
            .O(N__41067),
            .I(measured_delay_tr_10));
    LocalMux I__9124 (
            .O(N__41064),
            .I(measured_delay_tr_10));
    CascadeMux I__9123 (
            .O(N__41057),
            .I(N__41054));
    InMux I__9122 (
            .O(N__41054),
            .I(N__41051));
    LocalMux I__9121 (
            .O(N__41051),
            .I(N__41048));
    Odrv4 I__9120 (
            .O(N__41048),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__9119 (
            .O(N__41045),
            .I(N__41042));
    InMux I__9118 (
            .O(N__41042),
            .I(N__41039));
    LocalMux I__9117 (
            .O(N__41039),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__9116 (
            .O(N__41036),
            .I(N__41033));
    InMux I__9115 (
            .O(N__41033),
            .I(N__41030));
    LocalMux I__9114 (
            .O(N__41030),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__9113 (
            .O(N__41027),
            .I(N__41023));
    InMux I__9112 (
            .O(N__41026),
            .I(N__41020));
    LocalMux I__9111 (
            .O(N__41023),
            .I(N__41014));
    LocalMux I__9110 (
            .O(N__41020),
            .I(N__41014));
    InMux I__9109 (
            .O(N__41019),
            .I(N__41011));
    Odrv12 I__9108 (
            .O(N__41014),
            .I(measured_delay_tr_9));
    LocalMux I__9107 (
            .O(N__41011),
            .I(measured_delay_tr_9));
    CascadeMux I__9106 (
            .O(N__41006),
            .I(N__41003));
    InMux I__9105 (
            .O(N__41003),
            .I(N__41000));
    LocalMux I__9104 (
            .O(N__41000),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__9103 (
            .O(N__40997),
            .I(N__40994));
    InMux I__9102 (
            .O(N__40994),
            .I(N__40991));
    LocalMux I__9101 (
            .O(N__40991),
            .I(N__40988));
    Odrv4 I__9100 (
            .O(N__40988),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__9099 (
            .O(N__40985),
            .I(N__40982));
    InMux I__9098 (
            .O(N__40982),
            .I(N__40979));
    LocalMux I__9097 (
            .O(N__40979),
            .I(N__40976));
    Odrv4 I__9096 (
            .O(N__40976),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__9095 (
            .O(N__40973),
            .I(N__40970));
    InMux I__9094 (
            .O(N__40970),
            .I(N__40967));
    LocalMux I__9093 (
            .O(N__40967),
            .I(N__40964));
    Span4Mux_h I__9092 (
            .O(N__40964),
            .I(N__40961));
    Odrv4 I__9091 (
            .O(N__40961),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__9090 (
            .O(N__40958),
            .I(N__40955));
    InMux I__9089 (
            .O(N__40955),
            .I(N__40952));
    LocalMux I__9088 (
            .O(N__40952),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__9087 (
            .O(N__40949),
            .I(N__40946));
    InMux I__9086 (
            .O(N__40946),
            .I(N__40943));
    LocalMux I__9085 (
            .O(N__40943),
            .I(N__40940));
    Odrv4 I__9084 (
            .O(N__40940),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__9083 (
            .O(N__40937),
            .I(N__40934));
    InMux I__9082 (
            .O(N__40934),
            .I(N__40931));
    LocalMux I__9081 (
            .O(N__40931),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__9080 (
            .O(N__40928),
            .I(N__40925));
    InMux I__9079 (
            .O(N__40925),
            .I(N__40922));
    LocalMux I__9078 (
            .O(N__40922),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    InMux I__9077 (
            .O(N__40919),
            .I(N__40916));
    LocalMux I__9076 (
            .O(N__40916),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__9075 (
            .O(N__40913),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ));
    CascadeMux I__9074 (
            .O(N__40910),
            .I(N__40907));
    InMux I__9073 (
            .O(N__40907),
            .I(N__40904));
    LocalMux I__9072 (
            .O(N__40904),
            .I(N__40901));
    Odrv4 I__9071 (
            .O(N__40901),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    InMux I__9070 (
            .O(N__40898),
            .I(N__40895));
    LocalMux I__9069 (
            .O(N__40895),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__9068 (
            .O(N__40892),
            .I(N__40889));
    InMux I__9067 (
            .O(N__40889),
            .I(N__40886));
    LocalMux I__9066 (
            .O(N__40886),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__9065 (
            .O(N__40883),
            .I(N__40880));
    InMux I__9064 (
            .O(N__40880),
            .I(N__40877));
    LocalMux I__9063 (
            .O(N__40877),
            .I(N__40874));
    Odrv4 I__9062 (
            .O(N__40874),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__9061 (
            .O(N__40871),
            .I(N__40868));
    InMux I__9060 (
            .O(N__40868),
            .I(N__40865));
    LocalMux I__9059 (
            .O(N__40865),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__9058 (
            .O(N__40862),
            .I(N__40859));
    InMux I__9057 (
            .O(N__40859),
            .I(N__40856));
    LocalMux I__9056 (
            .O(N__40856),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    InMux I__9055 (
            .O(N__40853),
            .I(N__40839));
    InMux I__9054 (
            .O(N__40852),
            .I(N__40832));
    InMux I__9053 (
            .O(N__40851),
            .I(N__40832));
    InMux I__9052 (
            .O(N__40850),
            .I(N__40832));
    InMux I__9051 (
            .O(N__40849),
            .I(N__40822));
    InMux I__9050 (
            .O(N__40848),
            .I(N__40822));
    InMux I__9049 (
            .O(N__40847),
            .I(N__40822));
    InMux I__9048 (
            .O(N__40846),
            .I(N__40822));
    InMux I__9047 (
            .O(N__40845),
            .I(N__40817));
    InMux I__9046 (
            .O(N__40844),
            .I(N__40817));
    InMux I__9045 (
            .O(N__40843),
            .I(N__40812));
    InMux I__9044 (
            .O(N__40842),
            .I(N__40812));
    LocalMux I__9043 (
            .O(N__40839),
            .I(N__40809));
    LocalMux I__9042 (
            .O(N__40832),
            .I(N__40806));
    InMux I__9041 (
            .O(N__40831),
            .I(N__40803));
    LocalMux I__9040 (
            .O(N__40822),
            .I(N__40800));
    LocalMux I__9039 (
            .O(N__40817),
            .I(N__40795));
    LocalMux I__9038 (
            .O(N__40812),
            .I(N__40795));
    Span4Mux_v I__9037 (
            .O(N__40809),
            .I(N__40781));
    Span4Mux_h I__9036 (
            .O(N__40806),
            .I(N__40778));
    LocalMux I__9035 (
            .O(N__40803),
            .I(N__40775));
    Span4Mux_h I__9034 (
            .O(N__40800),
            .I(N__40772));
    Span4Mux_h I__9033 (
            .O(N__40795),
            .I(N__40769));
    InMux I__9032 (
            .O(N__40794),
            .I(N__40762));
    InMux I__9031 (
            .O(N__40793),
            .I(N__40762));
    InMux I__9030 (
            .O(N__40792),
            .I(N__40762));
    InMux I__9029 (
            .O(N__40791),
            .I(N__40745));
    InMux I__9028 (
            .O(N__40790),
            .I(N__40745));
    InMux I__9027 (
            .O(N__40789),
            .I(N__40745));
    InMux I__9026 (
            .O(N__40788),
            .I(N__40745));
    InMux I__9025 (
            .O(N__40787),
            .I(N__40745));
    InMux I__9024 (
            .O(N__40786),
            .I(N__40745));
    InMux I__9023 (
            .O(N__40785),
            .I(N__40745));
    InMux I__9022 (
            .O(N__40784),
            .I(N__40745));
    Odrv4 I__9021 (
            .O(N__40781),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__9020 (
            .O(N__40778),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv12 I__9019 (
            .O(N__40775),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__9018 (
            .O(N__40772),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__9017 (
            .O(N__40769),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__9016 (
            .O(N__40762),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__9015 (
            .O(N__40745),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    CascadeMux I__9014 (
            .O(N__40730),
            .I(N__40725));
    CascadeMux I__9013 (
            .O(N__40729),
            .I(N__40713));
    CascadeMux I__9012 (
            .O(N__40728),
            .I(N__40710));
    InMux I__9011 (
            .O(N__40725),
            .I(N__40706));
    InMux I__9010 (
            .O(N__40724),
            .I(N__40703));
    InMux I__9009 (
            .O(N__40723),
            .I(N__40688));
    InMux I__9008 (
            .O(N__40722),
            .I(N__40688));
    CascadeMux I__9007 (
            .O(N__40721),
            .I(N__40685));
    InMux I__9006 (
            .O(N__40720),
            .I(N__40672));
    InMux I__9005 (
            .O(N__40719),
            .I(N__40672));
    InMux I__9004 (
            .O(N__40718),
            .I(N__40672));
    InMux I__9003 (
            .O(N__40717),
            .I(N__40672));
    CascadeMux I__9002 (
            .O(N__40716),
            .I(N__40667));
    InMux I__9001 (
            .O(N__40713),
            .I(N__40659));
    InMux I__9000 (
            .O(N__40710),
            .I(N__40659));
    InMux I__8999 (
            .O(N__40709),
            .I(N__40659));
    LocalMux I__8998 (
            .O(N__40706),
            .I(N__40654));
    LocalMux I__8997 (
            .O(N__40703),
            .I(N__40654));
    InMux I__8996 (
            .O(N__40702),
            .I(N__40649));
    InMux I__8995 (
            .O(N__40701),
            .I(N__40632));
    InMux I__8994 (
            .O(N__40700),
            .I(N__40632));
    InMux I__8993 (
            .O(N__40699),
            .I(N__40632));
    InMux I__8992 (
            .O(N__40698),
            .I(N__40632));
    InMux I__8991 (
            .O(N__40697),
            .I(N__40632));
    InMux I__8990 (
            .O(N__40696),
            .I(N__40632));
    InMux I__8989 (
            .O(N__40695),
            .I(N__40632));
    InMux I__8988 (
            .O(N__40694),
            .I(N__40632));
    InMux I__8987 (
            .O(N__40693),
            .I(N__40629));
    LocalMux I__8986 (
            .O(N__40688),
            .I(N__40626));
    InMux I__8985 (
            .O(N__40685),
            .I(N__40615));
    InMux I__8984 (
            .O(N__40684),
            .I(N__40615));
    InMux I__8983 (
            .O(N__40683),
            .I(N__40615));
    InMux I__8982 (
            .O(N__40682),
            .I(N__40615));
    InMux I__8981 (
            .O(N__40681),
            .I(N__40615));
    LocalMux I__8980 (
            .O(N__40672),
            .I(N__40612));
    InMux I__8979 (
            .O(N__40671),
            .I(N__40603));
    InMux I__8978 (
            .O(N__40670),
            .I(N__40603));
    InMux I__8977 (
            .O(N__40667),
            .I(N__40603));
    InMux I__8976 (
            .O(N__40666),
            .I(N__40603));
    LocalMux I__8975 (
            .O(N__40659),
            .I(N__40600));
    Span4Mux_h I__8974 (
            .O(N__40654),
            .I(N__40597));
    InMux I__8973 (
            .O(N__40653),
            .I(N__40592));
    InMux I__8972 (
            .O(N__40652),
            .I(N__40592));
    LocalMux I__8971 (
            .O(N__40649),
            .I(N__40587));
    LocalMux I__8970 (
            .O(N__40632),
            .I(N__40587));
    LocalMux I__8969 (
            .O(N__40629),
            .I(N__40582));
    Span4Mux_h I__8968 (
            .O(N__40626),
            .I(N__40582));
    LocalMux I__8967 (
            .O(N__40615),
            .I(N__40577));
    Span4Mux_h I__8966 (
            .O(N__40612),
            .I(N__40577));
    LocalMux I__8965 (
            .O(N__40603),
            .I(N__40570));
    Span4Mux_h I__8964 (
            .O(N__40600),
            .I(N__40570));
    Span4Mux_h I__8963 (
            .O(N__40597),
            .I(N__40570));
    LocalMux I__8962 (
            .O(N__40592),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__8961 (
            .O(N__40587),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__8960 (
            .O(N__40582),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__8959 (
            .O(N__40577),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__8958 (
            .O(N__40570),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    CascadeMux I__8957 (
            .O(N__40559),
            .I(N__40555));
    CascadeMux I__8956 (
            .O(N__40558),
            .I(N__40548));
    InMux I__8955 (
            .O(N__40555),
            .I(N__40541));
    InMux I__8954 (
            .O(N__40554),
            .I(N__40541));
    CascadeMux I__8953 (
            .O(N__40553),
            .I(N__40538));
    CascadeMux I__8952 (
            .O(N__40552),
            .I(N__40526));
    CascadeMux I__8951 (
            .O(N__40551),
            .I(N__40521));
    InMux I__8950 (
            .O(N__40548),
            .I(N__40512));
    InMux I__8949 (
            .O(N__40547),
            .I(N__40512));
    InMux I__8948 (
            .O(N__40546),
            .I(N__40512));
    LocalMux I__8947 (
            .O(N__40541),
            .I(N__40506));
    InMux I__8946 (
            .O(N__40538),
            .I(N__40503));
    CascadeMux I__8945 (
            .O(N__40537),
            .I(N__40499));
    CascadeMux I__8944 (
            .O(N__40536),
            .I(N__40493));
    CascadeMux I__8943 (
            .O(N__40535),
            .I(N__40490));
    CascadeMux I__8942 (
            .O(N__40534),
            .I(N__40482));
    CascadeMux I__8941 (
            .O(N__40533),
            .I(N__40479));
    CascadeMux I__8940 (
            .O(N__40532),
            .I(N__40472));
    CascadeMux I__8939 (
            .O(N__40531),
            .I(N__40468));
    CascadeMux I__8938 (
            .O(N__40530),
            .I(N__40465));
    InMux I__8937 (
            .O(N__40529),
            .I(N__40458));
    InMux I__8936 (
            .O(N__40526),
            .I(N__40445));
    InMux I__8935 (
            .O(N__40525),
            .I(N__40445));
    InMux I__8934 (
            .O(N__40524),
            .I(N__40445));
    InMux I__8933 (
            .O(N__40521),
            .I(N__40445));
    InMux I__8932 (
            .O(N__40520),
            .I(N__40445));
    InMux I__8931 (
            .O(N__40519),
            .I(N__40445));
    LocalMux I__8930 (
            .O(N__40512),
            .I(N__40442));
    InMux I__8929 (
            .O(N__40511),
            .I(N__40437));
    InMux I__8928 (
            .O(N__40510),
            .I(N__40437));
    CascadeMux I__8927 (
            .O(N__40509),
            .I(N__40434));
    Sp12to4 I__8926 (
            .O(N__40506),
            .I(N__40429));
    LocalMux I__8925 (
            .O(N__40503),
            .I(N__40429));
    InMux I__8924 (
            .O(N__40502),
            .I(N__40418));
    InMux I__8923 (
            .O(N__40499),
            .I(N__40418));
    InMux I__8922 (
            .O(N__40498),
            .I(N__40418));
    InMux I__8921 (
            .O(N__40497),
            .I(N__40418));
    InMux I__8920 (
            .O(N__40496),
            .I(N__40418));
    InMux I__8919 (
            .O(N__40493),
            .I(N__40407));
    InMux I__8918 (
            .O(N__40490),
            .I(N__40407));
    InMux I__8917 (
            .O(N__40489),
            .I(N__40407));
    InMux I__8916 (
            .O(N__40488),
            .I(N__40407));
    InMux I__8915 (
            .O(N__40487),
            .I(N__40407));
    InMux I__8914 (
            .O(N__40486),
            .I(N__40390));
    InMux I__8913 (
            .O(N__40485),
            .I(N__40390));
    InMux I__8912 (
            .O(N__40482),
            .I(N__40390));
    InMux I__8911 (
            .O(N__40479),
            .I(N__40390));
    InMux I__8910 (
            .O(N__40478),
            .I(N__40390));
    InMux I__8909 (
            .O(N__40477),
            .I(N__40390));
    InMux I__8908 (
            .O(N__40476),
            .I(N__40390));
    InMux I__8907 (
            .O(N__40475),
            .I(N__40390));
    InMux I__8906 (
            .O(N__40472),
            .I(N__40385));
    InMux I__8905 (
            .O(N__40471),
            .I(N__40385));
    InMux I__8904 (
            .O(N__40468),
            .I(N__40374));
    InMux I__8903 (
            .O(N__40465),
            .I(N__40374));
    InMux I__8902 (
            .O(N__40464),
            .I(N__40374));
    InMux I__8901 (
            .O(N__40463),
            .I(N__40374));
    InMux I__8900 (
            .O(N__40462),
            .I(N__40374));
    InMux I__8899 (
            .O(N__40461),
            .I(N__40371));
    LocalMux I__8898 (
            .O(N__40458),
            .I(N__40362));
    LocalMux I__8897 (
            .O(N__40445),
            .I(N__40362));
    Span4Mux_v I__8896 (
            .O(N__40442),
            .I(N__40362));
    LocalMux I__8895 (
            .O(N__40437),
            .I(N__40362));
    InMux I__8894 (
            .O(N__40434),
            .I(N__40359));
    Span12Mux_s4_h I__8893 (
            .O(N__40429),
            .I(N__40355));
    LocalMux I__8892 (
            .O(N__40418),
            .I(N__40346));
    LocalMux I__8891 (
            .O(N__40407),
            .I(N__40346));
    LocalMux I__8890 (
            .O(N__40390),
            .I(N__40346));
    LocalMux I__8889 (
            .O(N__40385),
            .I(N__40346));
    LocalMux I__8888 (
            .O(N__40374),
            .I(N__40343));
    LocalMux I__8887 (
            .O(N__40371),
            .I(N__40340));
    Span4Mux_v I__8886 (
            .O(N__40362),
            .I(N__40335));
    LocalMux I__8885 (
            .O(N__40359),
            .I(N__40335));
    InMux I__8884 (
            .O(N__40358),
            .I(N__40332));
    Span12Mux_h I__8883 (
            .O(N__40355),
            .I(N__40329));
    Span4Mux_v I__8882 (
            .O(N__40346),
            .I(N__40326));
    Span4Mux_h I__8881 (
            .O(N__40343),
            .I(N__40323));
    Span4Mux_h I__8880 (
            .O(N__40340),
            .I(N__40318));
    Span4Mux_h I__8879 (
            .O(N__40335),
            .I(N__40318));
    LocalMux I__8878 (
            .O(N__40332),
            .I(measured_delay_hc_31));
    Odrv12 I__8877 (
            .O(N__40329),
            .I(measured_delay_hc_31));
    Odrv4 I__8876 (
            .O(N__40326),
            .I(measured_delay_hc_31));
    Odrv4 I__8875 (
            .O(N__40323),
            .I(measured_delay_hc_31));
    Odrv4 I__8874 (
            .O(N__40318),
            .I(measured_delay_hc_31));
    InMux I__8873 (
            .O(N__40307),
            .I(N__40304));
    LocalMux I__8872 (
            .O(N__40304),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__8871 (
            .O(N__40301),
            .I(N__40297));
    InMux I__8870 (
            .O(N__40300),
            .I(N__40294));
    LocalMux I__8869 (
            .O(N__40297),
            .I(N__40291));
    LocalMux I__8868 (
            .O(N__40294),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv12 I__8867 (
            .O(N__40291),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__8866 (
            .O(N__40286),
            .I(N__40283));
    LocalMux I__8865 (
            .O(N__40283),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__8864 (
            .O(N__40280),
            .I(N__40276));
    InMux I__8863 (
            .O(N__40279),
            .I(N__40273));
    LocalMux I__8862 (
            .O(N__40276),
            .I(N__40270));
    LocalMux I__8861 (
            .O(N__40273),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__8860 (
            .O(N__40270),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__8859 (
            .O(N__40265),
            .I(N__40262));
    LocalMux I__8858 (
            .O(N__40262),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__8857 (
            .O(N__40259),
            .I(N__40255));
    InMux I__8856 (
            .O(N__40258),
            .I(N__40252));
    LocalMux I__8855 (
            .O(N__40255),
            .I(N__40249));
    LocalMux I__8854 (
            .O(N__40252),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv12 I__8853 (
            .O(N__40249),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__8852 (
            .O(N__40244),
            .I(N__40220));
    InMux I__8851 (
            .O(N__40243),
            .I(N__40220));
    InMux I__8850 (
            .O(N__40242),
            .I(N__40220));
    InMux I__8849 (
            .O(N__40241),
            .I(N__40220));
    InMux I__8848 (
            .O(N__40240),
            .I(N__40203));
    InMux I__8847 (
            .O(N__40239),
            .I(N__40203));
    InMux I__8846 (
            .O(N__40238),
            .I(N__40203));
    InMux I__8845 (
            .O(N__40237),
            .I(N__40203));
    InMux I__8844 (
            .O(N__40236),
            .I(N__40203));
    InMux I__8843 (
            .O(N__40235),
            .I(N__40203));
    InMux I__8842 (
            .O(N__40234),
            .I(N__40203));
    InMux I__8841 (
            .O(N__40233),
            .I(N__40203));
    InMux I__8840 (
            .O(N__40232),
            .I(N__40194));
    InMux I__8839 (
            .O(N__40231),
            .I(N__40188));
    InMux I__8838 (
            .O(N__40230),
            .I(N__40188));
    CascadeMux I__8837 (
            .O(N__40229),
            .I(N__40185));
    LocalMux I__8836 (
            .O(N__40220),
            .I(N__40179));
    LocalMux I__8835 (
            .O(N__40203),
            .I(N__40179));
    InMux I__8834 (
            .O(N__40202),
            .I(N__40176));
    InMux I__8833 (
            .O(N__40201),
            .I(N__40165));
    InMux I__8832 (
            .O(N__40200),
            .I(N__40165));
    InMux I__8831 (
            .O(N__40199),
            .I(N__40165));
    InMux I__8830 (
            .O(N__40198),
            .I(N__40165));
    InMux I__8829 (
            .O(N__40197),
            .I(N__40165));
    LocalMux I__8828 (
            .O(N__40194),
            .I(N__40162));
    InMux I__8827 (
            .O(N__40193),
            .I(N__40159));
    LocalMux I__8826 (
            .O(N__40188),
            .I(N__40156));
    InMux I__8825 (
            .O(N__40185),
            .I(N__40151));
    InMux I__8824 (
            .O(N__40184),
            .I(N__40151));
    Span4Mux_h I__8823 (
            .O(N__40179),
            .I(N__40148));
    LocalMux I__8822 (
            .O(N__40176),
            .I(N__40145));
    LocalMux I__8821 (
            .O(N__40165),
            .I(N__40136));
    Span4Mux_v I__8820 (
            .O(N__40162),
            .I(N__40136));
    LocalMux I__8819 (
            .O(N__40159),
            .I(N__40136));
    Span4Mux_h I__8818 (
            .O(N__40156),
            .I(N__40136));
    LocalMux I__8817 (
            .O(N__40151),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8816 (
            .O(N__40148),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__8815 (
            .O(N__40145),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8814 (
            .O(N__40136),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__8813 (
            .O(N__40127),
            .I(N__40117));
    CascadeMux I__8812 (
            .O(N__40126),
            .I(N__40110));
    CascadeMux I__8811 (
            .O(N__40125),
            .I(N__40107));
    CascadeMux I__8810 (
            .O(N__40124),
            .I(N__40104));
    CascadeMux I__8809 (
            .O(N__40123),
            .I(N__40101));
    CascadeMux I__8808 (
            .O(N__40122),
            .I(N__40097));
    CascadeMux I__8807 (
            .O(N__40121),
            .I(N__40094));
    CascadeMux I__8806 (
            .O(N__40120),
            .I(N__40091));
    InMux I__8805 (
            .O(N__40117),
            .I(N__40087));
    InMux I__8804 (
            .O(N__40116),
            .I(N__40070));
    InMux I__8803 (
            .O(N__40115),
            .I(N__40070));
    InMux I__8802 (
            .O(N__40114),
            .I(N__40070));
    InMux I__8801 (
            .O(N__40113),
            .I(N__40070));
    InMux I__8800 (
            .O(N__40110),
            .I(N__40070));
    InMux I__8799 (
            .O(N__40107),
            .I(N__40070));
    InMux I__8798 (
            .O(N__40104),
            .I(N__40070));
    InMux I__8797 (
            .O(N__40101),
            .I(N__40070));
    CascadeMux I__8796 (
            .O(N__40100),
            .I(N__40067));
    InMux I__8795 (
            .O(N__40097),
            .I(N__40051));
    InMux I__8794 (
            .O(N__40094),
            .I(N__40051));
    InMux I__8793 (
            .O(N__40091),
            .I(N__40051));
    InMux I__8792 (
            .O(N__40090),
            .I(N__40051));
    LocalMux I__8791 (
            .O(N__40087),
            .I(N__40048));
    LocalMux I__8790 (
            .O(N__40070),
            .I(N__40045));
    InMux I__8789 (
            .O(N__40067),
            .I(N__40040));
    InMux I__8788 (
            .O(N__40066),
            .I(N__40040));
    InMux I__8787 (
            .O(N__40065),
            .I(N__40029));
    InMux I__8786 (
            .O(N__40064),
            .I(N__40029));
    InMux I__8785 (
            .O(N__40063),
            .I(N__40029));
    InMux I__8784 (
            .O(N__40062),
            .I(N__40029));
    InMux I__8783 (
            .O(N__40061),
            .I(N__40029));
    InMux I__8782 (
            .O(N__40060),
            .I(N__40026));
    LocalMux I__8781 (
            .O(N__40051),
            .I(N__40021));
    Span4Mux_v I__8780 (
            .O(N__40048),
            .I(N__40018));
    Span4Mux_h I__8779 (
            .O(N__40045),
            .I(N__40013));
    LocalMux I__8778 (
            .O(N__40040),
            .I(N__40013));
    LocalMux I__8777 (
            .O(N__40029),
            .I(N__40010));
    LocalMux I__8776 (
            .O(N__40026),
            .I(N__40007));
    InMux I__8775 (
            .O(N__40025),
            .I(N__40001));
    InMux I__8774 (
            .O(N__40024),
            .I(N__40001));
    Span4Mux_v I__8773 (
            .O(N__40021),
            .I(N__39996));
    Span4Mux_h I__8772 (
            .O(N__40018),
            .I(N__39996));
    Span4Mux_v I__8771 (
            .O(N__40013),
            .I(N__39991));
    Span4Mux_h I__8770 (
            .O(N__40010),
            .I(N__39991));
    Span4Mux_h I__8769 (
            .O(N__40007),
            .I(N__39988));
    InMux I__8768 (
            .O(N__40006),
            .I(N__39985));
    LocalMux I__8767 (
            .O(N__40001),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8766 (
            .O(N__39996),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8765 (
            .O(N__39991),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8764 (
            .O(N__39988),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__8763 (
            .O(N__39985),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__8762 (
            .O(N__39974),
            .I(N__39971));
    InMux I__8761 (
            .O(N__39971),
            .I(N__39968));
    LocalMux I__8760 (
            .O(N__39968),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__8759 (
            .O(N__39965),
            .I(N__39939));
    InMux I__8758 (
            .O(N__39964),
            .I(N__39939));
    InMux I__8757 (
            .O(N__39963),
            .I(N__39939));
    InMux I__8756 (
            .O(N__39962),
            .I(N__39939));
    CascadeMux I__8755 (
            .O(N__39961),
            .I(N__39933));
    CascadeMux I__8754 (
            .O(N__39960),
            .I(N__39930));
    CascadeMux I__8753 (
            .O(N__39959),
            .I(N__39927));
    InMux I__8752 (
            .O(N__39958),
            .I(N__39924));
    InMux I__8751 (
            .O(N__39957),
            .I(N__39920));
    InMux I__8750 (
            .O(N__39956),
            .I(N__39917));
    InMux I__8749 (
            .O(N__39955),
            .I(N__39898));
    InMux I__8748 (
            .O(N__39954),
            .I(N__39898));
    InMux I__8747 (
            .O(N__39953),
            .I(N__39898));
    InMux I__8746 (
            .O(N__39952),
            .I(N__39898));
    InMux I__8745 (
            .O(N__39951),
            .I(N__39898));
    InMux I__8744 (
            .O(N__39950),
            .I(N__39898));
    InMux I__8743 (
            .O(N__39949),
            .I(N__39898));
    InMux I__8742 (
            .O(N__39948),
            .I(N__39898));
    LocalMux I__8741 (
            .O(N__39939),
            .I(N__39895));
    InMux I__8740 (
            .O(N__39938),
            .I(N__39892));
    InMux I__8739 (
            .O(N__39937),
            .I(N__39881));
    InMux I__8738 (
            .O(N__39936),
            .I(N__39881));
    InMux I__8737 (
            .O(N__39933),
            .I(N__39881));
    InMux I__8736 (
            .O(N__39930),
            .I(N__39881));
    InMux I__8735 (
            .O(N__39927),
            .I(N__39881));
    LocalMux I__8734 (
            .O(N__39924),
            .I(N__39878));
    InMux I__8733 (
            .O(N__39923),
            .I(N__39875));
    LocalMux I__8732 (
            .O(N__39920),
            .I(N__39870));
    LocalMux I__8731 (
            .O(N__39917),
            .I(N__39870));
    InMux I__8730 (
            .O(N__39916),
            .I(N__39865));
    InMux I__8729 (
            .O(N__39915),
            .I(N__39865));
    LocalMux I__8728 (
            .O(N__39898),
            .I(N__39862));
    Span4Mux_h I__8727 (
            .O(N__39895),
            .I(N__39859));
    LocalMux I__8726 (
            .O(N__39892),
            .I(N__39856));
    LocalMux I__8725 (
            .O(N__39881),
            .I(N__39847));
    Span4Mux_v I__8724 (
            .O(N__39878),
            .I(N__39847));
    LocalMux I__8723 (
            .O(N__39875),
            .I(N__39847));
    Span4Mux_h I__8722 (
            .O(N__39870),
            .I(N__39847));
    LocalMux I__8721 (
            .O(N__39865),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__8720 (
            .O(N__39862),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__8719 (
            .O(N__39859),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv12 I__8718 (
            .O(N__39856),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__8717 (
            .O(N__39847),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__8716 (
            .O(N__39836),
            .I(N__39833));
    LocalMux I__8715 (
            .O(N__39833),
            .I(N__39829));
    InMux I__8714 (
            .O(N__39832),
            .I(N__39826));
    Span4Mux_h I__8713 (
            .O(N__39829),
            .I(N__39823));
    LocalMux I__8712 (
            .O(N__39826),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__8711 (
            .O(N__39823),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CEMux I__8710 (
            .O(N__39818),
            .I(N__39814));
    CEMux I__8709 (
            .O(N__39817),
            .I(N__39811));
    LocalMux I__8708 (
            .O(N__39814),
            .I(N__39808));
    LocalMux I__8707 (
            .O(N__39811),
            .I(N__39805));
    Span4Mux_v I__8706 (
            .O(N__39808),
            .I(N__39802));
    Span4Mux_h I__8705 (
            .O(N__39805),
            .I(N__39798));
    Span4Mux_h I__8704 (
            .O(N__39802),
            .I(N__39795));
    CEMux I__8703 (
            .O(N__39801),
            .I(N__39792));
    Span4Mux_h I__8702 (
            .O(N__39798),
            .I(N__39789));
    Sp12to4 I__8701 (
            .O(N__39795),
            .I(N__39784));
    LocalMux I__8700 (
            .O(N__39792),
            .I(N__39784));
    Odrv4 I__8699 (
            .O(N__39789),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv12 I__8698 (
            .O(N__39784),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__8697 (
            .O(N__39779),
            .I(N__39776));
    LocalMux I__8696 (
            .O(N__39776),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_0 ));
    CascadeMux I__8695 (
            .O(N__39773),
            .I(\delay_measurement_inst.delay_hc_reg3lto30_2_cascade_ ));
    CascadeMux I__8694 (
            .O(N__39770),
            .I(\delay_measurement_inst.delay_hc_reg3_cascade_ ));
    InMux I__8693 (
            .O(N__39767),
            .I(N__39763));
    InMux I__8692 (
            .O(N__39766),
            .I(N__39760));
    LocalMux I__8691 (
            .O(N__39763),
            .I(N__39755));
    LocalMux I__8690 (
            .O(N__39760),
            .I(N__39752));
    InMux I__8689 (
            .O(N__39759),
            .I(N__39749));
    InMux I__8688 (
            .O(N__39758),
            .I(N__39746));
    Span12Mux_v I__8687 (
            .O(N__39755),
            .I(N__39743));
    Span4Mux_h I__8686 (
            .O(N__39752),
            .I(N__39740));
    LocalMux I__8685 (
            .O(N__39749),
            .I(N__39737));
    LocalMux I__8684 (
            .O(N__39746),
            .I(measured_delay_hc_4));
    Odrv12 I__8683 (
            .O(N__39743),
            .I(measured_delay_hc_4));
    Odrv4 I__8682 (
            .O(N__39740),
            .I(measured_delay_hc_4));
    Odrv4 I__8681 (
            .O(N__39737),
            .I(measured_delay_hc_4));
    CascadeMux I__8680 (
            .O(N__39728),
            .I(N__39725));
    InMux I__8679 (
            .O(N__39725),
            .I(N__39719));
    InMux I__8678 (
            .O(N__39724),
            .I(N__39716));
    CascadeMux I__8677 (
            .O(N__39723),
            .I(N__39713));
    InMux I__8676 (
            .O(N__39722),
            .I(N__39709));
    LocalMux I__8675 (
            .O(N__39719),
            .I(N__39704));
    LocalMux I__8674 (
            .O(N__39716),
            .I(N__39704));
    InMux I__8673 (
            .O(N__39713),
            .I(N__39701));
    CascadeMux I__8672 (
            .O(N__39712),
            .I(N__39698));
    LocalMux I__8671 (
            .O(N__39709),
            .I(N__39695));
    Span4Mux_v I__8670 (
            .O(N__39704),
            .I(N__39690));
    LocalMux I__8669 (
            .O(N__39701),
            .I(N__39690));
    InMux I__8668 (
            .O(N__39698),
            .I(N__39687));
    Span4Mux_h I__8667 (
            .O(N__39695),
            .I(N__39682));
    Span4Mux_h I__8666 (
            .O(N__39690),
            .I(N__39682));
    LocalMux I__8665 (
            .O(N__39687),
            .I(measured_delay_hc_14));
    Odrv4 I__8664 (
            .O(N__39682),
            .I(measured_delay_hc_14));
    InMux I__8663 (
            .O(N__39677),
            .I(N__39674));
    LocalMux I__8662 (
            .O(N__39674),
            .I(N__39670));
    InMux I__8661 (
            .O(N__39673),
            .I(N__39667));
    Span4Mux_v I__8660 (
            .O(N__39670),
            .I(N__39664));
    LocalMux I__8659 (
            .O(N__39667),
            .I(measured_delay_hc_24));
    Odrv4 I__8658 (
            .O(N__39664),
            .I(measured_delay_hc_24));
    InMux I__8657 (
            .O(N__39659),
            .I(N__39656));
    LocalMux I__8656 (
            .O(N__39656),
            .I(N__39652));
    InMux I__8655 (
            .O(N__39655),
            .I(N__39649));
    Span4Mux_h I__8654 (
            .O(N__39652),
            .I(N__39646));
    LocalMux I__8653 (
            .O(N__39649),
            .I(measured_delay_hc_25));
    Odrv4 I__8652 (
            .O(N__39646),
            .I(measured_delay_hc_25));
    CascadeMux I__8651 (
            .O(N__39641),
            .I(N__39638));
    InMux I__8650 (
            .O(N__39638),
            .I(N__39635));
    LocalMux I__8649 (
            .O(N__39635),
            .I(N__39631));
    InMux I__8648 (
            .O(N__39634),
            .I(N__39628));
    Span4Mux_h I__8647 (
            .O(N__39631),
            .I(N__39625));
    LocalMux I__8646 (
            .O(N__39628),
            .I(measured_delay_hc_26));
    Odrv4 I__8645 (
            .O(N__39625),
            .I(measured_delay_hc_26));
    InMux I__8644 (
            .O(N__39620),
            .I(N__39616));
    InMux I__8643 (
            .O(N__39619),
            .I(N__39613));
    LocalMux I__8642 (
            .O(N__39616),
            .I(measured_delay_hc_28));
    LocalMux I__8641 (
            .O(N__39613),
            .I(measured_delay_hc_28));
    InMux I__8640 (
            .O(N__39608),
            .I(N__39604));
    InMux I__8639 (
            .O(N__39607),
            .I(N__39601));
    LocalMux I__8638 (
            .O(N__39604),
            .I(measured_delay_hc_30));
    LocalMux I__8637 (
            .O(N__39601),
            .I(measured_delay_hc_30));
    InMux I__8636 (
            .O(N__39596),
            .I(N__39593));
    LocalMux I__8635 (
            .O(N__39593),
            .I(N__39588));
    InMux I__8634 (
            .O(N__39592),
            .I(N__39585));
    InMux I__8633 (
            .O(N__39591),
            .I(N__39582));
    Span12Mux_v I__8632 (
            .O(N__39588),
            .I(N__39578));
    LocalMux I__8631 (
            .O(N__39585),
            .I(N__39575));
    LocalMux I__8630 (
            .O(N__39582),
            .I(N__39572));
    InMux I__8629 (
            .O(N__39581),
            .I(N__39569));
    Span12Mux_h I__8628 (
            .O(N__39578),
            .I(N__39566));
    Span4Mux_h I__8627 (
            .O(N__39575),
            .I(N__39563));
    Span4Mux_h I__8626 (
            .O(N__39572),
            .I(N__39560));
    LocalMux I__8625 (
            .O(N__39569),
            .I(measured_delay_hc_0));
    Odrv12 I__8624 (
            .O(N__39566),
            .I(measured_delay_hc_0));
    Odrv4 I__8623 (
            .O(N__39563),
            .I(measured_delay_hc_0));
    Odrv4 I__8622 (
            .O(N__39560),
            .I(measured_delay_hc_0));
    InMux I__8621 (
            .O(N__39551),
            .I(N__39527));
    InMux I__8620 (
            .O(N__39550),
            .I(N__39527));
    InMux I__8619 (
            .O(N__39549),
            .I(N__39527));
    InMux I__8618 (
            .O(N__39548),
            .I(N__39527));
    InMux I__8617 (
            .O(N__39547),
            .I(N__39518));
    InMux I__8616 (
            .O(N__39546),
            .I(N__39518));
    InMux I__8615 (
            .O(N__39545),
            .I(N__39518));
    InMux I__8614 (
            .O(N__39544),
            .I(N__39518));
    InMux I__8613 (
            .O(N__39543),
            .I(N__39495));
    InMux I__8612 (
            .O(N__39542),
            .I(N__39495));
    InMux I__8611 (
            .O(N__39541),
            .I(N__39495));
    InMux I__8610 (
            .O(N__39540),
            .I(N__39495));
    InMux I__8609 (
            .O(N__39539),
            .I(N__39486));
    InMux I__8608 (
            .O(N__39538),
            .I(N__39486));
    InMux I__8607 (
            .O(N__39537),
            .I(N__39486));
    InMux I__8606 (
            .O(N__39536),
            .I(N__39486));
    LocalMux I__8605 (
            .O(N__39527),
            .I(N__39481));
    LocalMux I__8604 (
            .O(N__39518),
            .I(N__39481));
    InMux I__8603 (
            .O(N__39517),
            .I(N__39472));
    InMux I__8602 (
            .O(N__39516),
            .I(N__39472));
    InMux I__8601 (
            .O(N__39515),
            .I(N__39472));
    InMux I__8600 (
            .O(N__39514),
            .I(N__39472));
    InMux I__8599 (
            .O(N__39513),
            .I(N__39467));
    InMux I__8598 (
            .O(N__39512),
            .I(N__39467));
    InMux I__8597 (
            .O(N__39511),
            .I(N__39458));
    InMux I__8596 (
            .O(N__39510),
            .I(N__39458));
    InMux I__8595 (
            .O(N__39509),
            .I(N__39458));
    InMux I__8594 (
            .O(N__39508),
            .I(N__39458));
    InMux I__8593 (
            .O(N__39507),
            .I(N__39449));
    InMux I__8592 (
            .O(N__39506),
            .I(N__39449));
    InMux I__8591 (
            .O(N__39505),
            .I(N__39449));
    InMux I__8590 (
            .O(N__39504),
            .I(N__39449));
    LocalMux I__8589 (
            .O(N__39495),
            .I(N__39444));
    LocalMux I__8588 (
            .O(N__39486),
            .I(N__39444));
    Sp12to4 I__8587 (
            .O(N__39481),
            .I(N__39435));
    LocalMux I__8586 (
            .O(N__39472),
            .I(N__39435));
    LocalMux I__8585 (
            .O(N__39467),
            .I(N__39435));
    LocalMux I__8584 (
            .O(N__39458),
            .I(N__39435));
    LocalMux I__8583 (
            .O(N__39449),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8582 (
            .O(N__39444),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv12 I__8581 (
            .O(N__39435),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__8580 (
            .O(N__39428),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CEMux I__8579 (
            .O(N__39425),
            .I(N__39420));
    CEMux I__8578 (
            .O(N__39424),
            .I(N__39417));
    CEMux I__8577 (
            .O(N__39423),
            .I(N__39414));
    LocalMux I__8576 (
            .O(N__39420),
            .I(N__39411));
    LocalMux I__8575 (
            .O(N__39417),
            .I(N__39406));
    LocalMux I__8574 (
            .O(N__39414),
            .I(N__39406));
    Span4Mux_v I__8573 (
            .O(N__39411),
            .I(N__39402));
    Span4Mux_v I__8572 (
            .O(N__39406),
            .I(N__39399));
    CEMux I__8571 (
            .O(N__39405),
            .I(N__39396));
    Odrv4 I__8570 (
            .O(N__39402),
            .I(\delay_measurement_inst.delay_hc_timer.N_336_i ));
    Odrv4 I__8569 (
            .O(N__39399),
            .I(\delay_measurement_inst.delay_hc_timer.N_336_i ));
    LocalMux I__8568 (
            .O(N__39396),
            .I(\delay_measurement_inst.delay_hc_timer.N_336_i ));
    CascadeMux I__8567 (
            .O(N__39389),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_ ));
    CascadeMux I__8566 (
            .O(N__39386),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_0_cascade_ ));
    CascadeMux I__8565 (
            .O(N__39383),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_cascade_ ));
    CascadeMux I__8564 (
            .O(N__39380),
            .I(N__39377));
    InMux I__8563 (
            .O(N__39377),
            .I(N__39374));
    LocalMux I__8562 (
            .O(N__39374),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ));
    InMux I__8561 (
            .O(N__39371),
            .I(N__39368));
    LocalMux I__8560 (
            .O(N__39368),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4 ));
    InMux I__8559 (
            .O(N__39365),
            .I(N__39361));
    InMux I__8558 (
            .O(N__39364),
            .I(N__39358));
    LocalMux I__8557 (
            .O(N__39361),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ));
    LocalMux I__8556 (
            .O(N__39358),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ));
    CascadeMux I__8555 (
            .O(N__39353),
            .I(N__39349));
    InMux I__8554 (
            .O(N__39352),
            .I(N__39346));
    InMux I__8553 (
            .O(N__39349),
            .I(N__39343));
    LocalMux I__8552 (
            .O(N__39346),
            .I(N__39340));
    LocalMux I__8551 (
            .O(N__39343),
            .I(N__39337));
    Span4Mux_v I__8550 (
            .O(N__39340),
            .I(N__39332));
    Span4Mux_h I__8549 (
            .O(N__39337),
            .I(N__39332));
    Span4Mux_h I__8548 (
            .O(N__39332),
            .I(N__39329));
    Span4Mux_h I__8547 (
            .O(N__39329),
            .I(N__39326));
    Odrv4 I__8546 (
            .O(N__39326),
            .I(\delay_measurement_inst.delay_hc_reg3lto30_2 ));
    InMux I__8545 (
            .O(N__39323),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__8544 (
            .O(N__39320),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__8543 (
            .O(N__39317),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__8542 (
            .O(N__39314),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__8541 (
            .O(N__39311),
            .I(bfn_16_10_0_));
    InMux I__8540 (
            .O(N__39308),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__8539 (
            .O(N__39305),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__8538 (
            .O(N__39302),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__8537 (
            .O(N__39299),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__8536 (
            .O(N__39296),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__8535 (
            .O(N__39293),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__8534 (
            .O(N__39290),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__8533 (
            .O(N__39287),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__8532 (
            .O(N__39284),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__8531 (
            .O(N__39281),
            .I(bfn_16_9_0_));
    InMux I__8530 (
            .O(N__39278),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__8529 (
            .O(N__39275),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__8528 (
            .O(N__39272),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__8527 (
            .O(N__39269),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__8526 (
            .O(N__39266),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__8525 (
            .O(N__39263),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__8524 (
            .O(N__39260),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__8523 (
            .O(N__39257),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__8522 (
            .O(N__39254),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__8521 (
            .O(N__39251),
            .I(bfn_16_8_0_));
    InMux I__8520 (
            .O(N__39248),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__8519 (
            .O(N__39245),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__8518 (
            .O(N__39242),
            .I(N__39238));
    InMux I__8517 (
            .O(N__39241),
            .I(N__39235));
    LocalMux I__8516 (
            .O(N__39238),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__8515 (
            .O(N__39235),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__8514 (
            .O(N__39230),
            .I(N__39227));
    LocalMux I__8513 (
            .O(N__39227),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__8512 (
            .O(N__39224),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__8511 (
            .O(N__39221),
            .I(N__39216));
    InMux I__8510 (
            .O(N__39220),
            .I(N__39213));
    InMux I__8509 (
            .O(N__39219),
            .I(N__39210));
    LocalMux I__8508 (
            .O(N__39216),
            .I(N__39207));
    LocalMux I__8507 (
            .O(N__39213),
            .I(N__39202));
    LocalMux I__8506 (
            .O(N__39210),
            .I(N__39198));
    Sp12to4 I__8505 (
            .O(N__39207),
            .I(N__39195));
    InMux I__8504 (
            .O(N__39206),
            .I(N__39190));
    InMux I__8503 (
            .O(N__39205),
            .I(N__39190));
    Span4Mux_h I__8502 (
            .O(N__39202),
            .I(N__39187));
    InMux I__8501 (
            .O(N__39201),
            .I(N__39184));
    Span12Mux_h I__8500 (
            .O(N__39198),
            .I(N__39179));
    Span12Mux_v I__8499 (
            .O(N__39195),
            .I(N__39179));
    LocalMux I__8498 (
            .O(N__39190),
            .I(N__39176));
    Odrv4 I__8497 (
            .O(N__39187),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__8496 (
            .O(N__39184),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__8495 (
            .O(N__39179),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__8494 (
            .O(N__39176),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__8493 (
            .O(N__39167),
            .I(N__39164));
    InMux I__8492 (
            .O(N__39164),
            .I(N__39161));
    LocalMux I__8491 (
            .O(N__39161),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__8490 (
            .O(N__39158),
            .I(N__39155));
    InMux I__8489 (
            .O(N__39155),
            .I(N__39152));
    LocalMux I__8488 (
            .O(N__39152),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__8487 (
            .O(N__39149),
            .I(N__39146));
    InMux I__8486 (
            .O(N__39146),
            .I(N__39143));
    LocalMux I__8485 (
            .O(N__39143),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__8484 (
            .O(N__39140),
            .I(N__39136));
    InMux I__8483 (
            .O(N__39139),
            .I(N__39133));
    LocalMux I__8482 (
            .O(N__39136),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__8481 (
            .O(N__39133),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__8480 (
            .O(N__39128),
            .I(N__39123));
    InMux I__8479 (
            .O(N__39127),
            .I(N__39120));
    InMux I__8478 (
            .O(N__39126),
            .I(N__39117));
    LocalMux I__8477 (
            .O(N__39123),
            .I(N__39114));
    LocalMux I__8476 (
            .O(N__39120),
            .I(N__39111));
    LocalMux I__8475 (
            .O(N__39117),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__8474 (
            .O(N__39114),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__8473 (
            .O(N__39111),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__8472 (
            .O(N__39104),
            .I(N__39098));
    InMux I__8471 (
            .O(N__39103),
            .I(N__39095));
    InMux I__8470 (
            .O(N__39102),
            .I(N__39090));
    InMux I__8469 (
            .O(N__39101),
            .I(N__39090));
    LocalMux I__8468 (
            .O(N__39098),
            .I(N__39087));
    LocalMux I__8467 (
            .O(N__39095),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__8466 (
            .O(N__39090),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__8465 (
            .O(N__39087),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__8464 (
            .O(N__39080),
            .I(bfn_16_7_0_));
    InMux I__8463 (
            .O(N__39077),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__8462 (
            .O(N__39074),
            .I(N__39070));
    InMux I__8461 (
            .O(N__39073),
            .I(N__39067));
    LocalMux I__8460 (
            .O(N__39070),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__8459 (
            .O(N__39067),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8458 (
            .O(N__39062),
            .I(N__39059));
    LocalMux I__8457 (
            .O(N__39059),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__8456 (
            .O(N__39056),
            .I(N__39052));
    InMux I__8455 (
            .O(N__39055),
            .I(N__39049));
    LocalMux I__8454 (
            .O(N__39052),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__8453 (
            .O(N__39049),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8452 (
            .O(N__39044),
            .I(N__39041));
    LocalMux I__8451 (
            .O(N__39041),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__8450 (
            .O(N__39038),
            .I(N__39034));
    InMux I__8449 (
            .O(N__39037),
            .I(N__39031));
    LocalMux I__8448 (
            .O(N__39034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__8447 (
            .O(N__39031),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8446 (
            .O(N__39026),
            .I(N__39023));
    LocalMux I__8445 (
            .O(N__39023),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__8444 (
            .O(N__39020),
            .I(N__39016));
    InMux I__8443 (
            .O(N__39019),
            .I(N__39013));
    LocalMux I__8442 (
            .O(N__39016),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__8441 (
            .O(N__39013),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8440 (
            .O(N__39008),
            .I(N__39005));
    LocalMux I__8439 (
            .O(N__39005),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__8438 (
            .O(N__39002),
            .I(N__38998));
    InMux I__8437 (
            .O(N__39001),
            .I(N__38995));
    LocalMux I__8436 (
            .O(N__38998),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__8435 (
            .O(N__38995),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__8434 (
            .O(N__38990),
            .I(N__38987));
    InMux I__8433 (
            .O(N__38987),
            .I(N__38984));
    LocalMux I__8432 (
            .O(N__38984),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__8431 (
            .O(N__38981),
            .I(N__38978));
    InMux I__8430 (
            .O(N__38978),
            .I(N__38975));
    LocalMux I__8429 (
            .O(N__38975),
            .I(N__38972));
    Odrv4 I__8428 (
            .O(N__38972),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__8427 (
            .O(N__38969),
            .I(N__38965));
    InMux I__8426 (
            .O(N__38968),
            .I(N__38962));
    LocalMux I__8425 (
            .O(N__38965),
            .I(N__38959));
    LocalMux I__8424 (
            .O(N__38962),
            .I(N__38954));
    Span4Mux_h I__8423 (
            .O(N__38959),
            .I(N__38954));
    Odrv4 I__8422 (
            .O(N__38954),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__8421 (
            .O(N__38951),
            .I(N__38948));
    LocalMux I__8420 (
            .O(N__38948),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    InMux I__8419 (
            .O(N__38945),
            .I(N__38941));
    InMux I__8418 (
            .O(N__38944),
            .I(N__38938));
    LocalMux I__8417 (
            .O(N__38941),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__8416 (
            .O(N__38938),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8415 (
            .O(N__38933),
            .I(N__38930));
    LocalMux I__8414 (
            .O(N__38930),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__8413 (
            .O(N__38927),
            .I(N__38923));
    InMux I__8412 (
            .O(N__38926),
            .I(N__38920));
    LocalMux I__8411 (
            .O(N__38923),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__8410 (
            .O(N__38920),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__8409 (
            .O(N__38915),
            .I(N__38912));
    LocalMux I__8408 (
            .O(N__38912),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__8407 (
            .O(N__38909),
            .I(N__38905));
    InMux I__8406 (
            .O(N__38908),
            .I(N__38902));
    LocalMux I__8405 (
            .O(N__38905),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__8404 (
            .O(N__38902),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8403 (
            .O(N__38897),
            .I(N__38894));
    LocalMux I__8402 (
            .O(N__38894),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__8401 (
            .O(N__38891),
            .I(N__38887));
    InMux I__8400 (
            .O(N__38890),
            .I(N__38884));
    LocalMux I__8399 (
            .O(N__38887),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__8398 (
            .O(N__38884),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8397 (
            .O(N__38879),
            .I(N__38876));
    LocalMux I__8396 (
            .O(N__38876),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__8395 (
            .O(N__38873),
            .I(N__38869));
    InMux I__8394 (
            .O(N__38872),
            .I(N__38866));
    LocalMux I__8393 (
            .O(N__38869),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__8392 (
            .O(N__38866),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__8391 (
            .O(N__38861),
            .I(N__38858));
    InMux I__8390 (
            .O(N__38858),
            .I(N__38855));
    LocalMux I__8389 (
            .O(N__38855),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__8388 (
            .O(N__38852),
            .I(N__38848));
    InMux I__8387 (
            .O(N__38851),
            .I(N__38845));
    LocalMux I__8386 (
            .O(N__38848),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__8385 (
            .O(N__38845),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8384 (
            .O(N__38840),
            .I(N__38837));
    LocalMux I__8383 (
            .O(N__38837),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__8382 (
            .O(N__38834),
            .I(N__38830));
    InMux I__8381 (
            .O(N__38833),
            .I(N__38827));
    LocalMux I__8380 (
            .O(N__38830),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__8379 (
            .O(N__38827),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8378 (
            .O(N__38822),
            .I(N__38819));
    LocalMux I__8377 (
            .O(N__38819),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__8376 (
            .O(N__38816),
            .I(N__38813));
    InMux I__8375 (
            .O(N__38813),
            .I(N__38809));
    InMux I__8374 (
            .O(N__38812),
            .I(N__38806));
    LocalMux I__8373 (
            .O(N__38809),
            .I(N__38803));
    LocalMux I__8372 (
            .O(N__38806),
            .I(N__38800));
    Odrv4 I__8371 (
            .O(N__38803),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__8370 (
            .O(N__38800),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8369 (
            .O(N__38795),
            .I(N__38792));
    LocalMux I__8368 (
            .O(N__38792),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__8367 (
            .O(N__38789),
            .I(N__38785));
    InMux I__8366 (
            .O(N__38788),
            .I(N__38782));
    LocalMux I__8365 (
            .O(N__38785),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__8364 (
            .O(N__38782),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8363 (
            .O(N__38777),
            .I(N__38774));
    LocalMux I__8362 (
            .O(N__38774),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__8361 (
            .O(N__38771),
            .I(N__38768));
    LocalMux I__8360 (
            .O(N__38768),
            .I(N__38764));
    InMux I__8359 (
            .O(N__38767),
            .I(N__38761));
    Span4Mux_h I__8358 (
            .O(N__38764),
            .I(N__38758));
    LocalMux I__8357 (
            .O(N__38761),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__8356 (
            .O(N__38758),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8355 (
            .O(N__38753),
            .I(N__38750));
    LocalMux I__8354 (
            .O(N__38750),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    InMux I__8353 (
            .O(N__38747),
            .I(N__38744));
    LocalMux I__8352 (
            .O(N__38744),
            .I(N__38740));
    InMux I__8351 (
            .O(N__38743),
            .I(N__38737));
    Span4Mux_h I__8350 (
            .O(N__38740),
            .I(N__38734));
    LocalMux I__8349 (
            .O(N__38737),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__8348 (
            .O(N__38734),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__8347 (
            .O(N__38729),
            .I(N__38726));
    LocalMux I__8346 (
            .O(N__38726),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    InMux I__8345 (
            .O(N__38723),
            .I(N__38719));
    InMux I__8344 (
            .O(N__38722),
            .I(N__38716));
    LocalMux I__8343 (
            .O(N__38719),
            .I(N__38713));
    LocalMux I__8342 (
            .O(N__38716),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__8341 (
            .O(N__38713),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__8340 (
            .O(N__38708),
            .I(N__38705));
    LocalMux I__8339 (
            .O(N__38705),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__8338 (
            .O(N__38702),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__8337 (
            .O(N__38699),
            .I(N__38692));
    InMux I__8336 (
            .O(N__38698),
            .I(N__38692));
    InMux I__8335 (
            .O(N__38697),
            .I(N__38689));
    LocalMux I__8334 (
            .O(N__38692),
            .I(N__38686));
    LocalMux I__8333 (
            .O(N__38689),
            .I(N__38683));
    Span4Mux_v I__8332 (
            .O(N__38686),
            .I(N__38677));
    Span4Mux_h I__8331 (
            .O(N__38683),
            .I(N__38674));
    InMux I__8330 (
            .O(N__38682),
            .I(N__38671));
    InMux I__8329 (
            .O(N__38681),
            .I(N__38668));
    InMux I__8328 (
            .O(N__38680),
            .I(N__38665));
    Span4Mux_v I__8327 (
            .O(N__38677),
            .I(N__38662));
    Span4Mux_v I__8326 (
            .O(N__38674),
            .I(N__38659));
    LocalMux I__8325 (
            .O(N__38671),
            .I(N__38656));
    LocalMux I__8324 (
            .O(N__38668),
            .I(N__38651));
    LocalMux I__8323 (
            .O(N__38665),
            .I(N__38651));
    Odrv4 I__8322 (
            .O(N__38662),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__8321 (
            .O(N__38659),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__8320 (
            .O(N__38656),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__8319 (
            .O(N__38651),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__8318 (
            .O(N__38642),
            .I(N__38639));
    InMux I__8317 (
            .O(N__38639),
            .I(N__38636));
    LocalMux I__8316 (
            .O(N__38636),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__8315 (
            .O(N__38633),
            .I(N__38630));
    InMux I__8314 (
            .O(N__38630),
            .I(N__38627));
    LocalMux I__8313 (
            .O(N__38627),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    InMux I__8312 (
            .O(N__38624),
            .I(N__38621));
    LocalMux I__8311 (
            .O(N__38621),
            .I(N__38617));
    CascadeMux I__8310 (
            .O(N__38620),
            .I(N__38614));
    Span12Mux_v I__8309 (
            .O(N__38617),
            .I(N__38610));
    InMux I__8308 (
            .O(N__38614),
            .I(N__38607));
    InMux I__8307 (
            .O(N__38613),
            .I(N__38604));
    Odrv12 I__8306 (
            .O(N__38610),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8305 (
            .O(N__38607),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8304 (
            .O(N__38604),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8303 (
            .O(N__38597),
            .I(N__38594));
    LocalMux I__8302 (
            .O(N__38594),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__8301 (
            .O(N__38591),
            .I(N__38587));
    InMux I__8300 (
            .O(N__38590),
            .I(N__38584));
    LocalMux I__8299 (
            .O(N__38587),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__8298 (
            .O(N__38584),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__8297 (
            .O(N__38579),
            .I(N__38576));
    InMux I__8296 (
            .O(N__38576),
            .I(N__38573));
    LocalMux I__8295 (
            .O(N__38573),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__8294 (
            .O(N__38570),
            .I(N__38567));
    InMux I__8293 (
            .O(N__38567),
            .I(N__38563));
    InMux I__8292 (
            .O(N__38566),
            .I(N__38560));
    LocalMux I__8291 (
            .O(N__38563),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__8290 (
            .O(N__38560),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8289 (
            .O(N__38555),
            .I(N__38552));
    LocalMux I__8288 (
            .O(N__38552),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__8287 (
            .O(N__38549),
            .I(N__38545));
    InMux I__8286 (
            .O(N__38548),
            .I(N__38542));
    LocalMux I__8285 (
            .O(N__38545),
            .I(N__38539));
    LocalMux I__8284 (
            .O(N__38542),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__8283 (
            .O(N__38539),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8282 (
            .O(N__38534),
            .I(N__38531));
    LocalMux I__8281 (
            .O(N__38531),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    InMux I__8280 (
            .O(N__38528),
            .I(N__38524));
    InMux I__8279 (
            .O(N__38527),
            .I(N__38521));
    LocalMux I__8278 (
            .O(N__38524),
            .I(N__38518));
    LocalMux I__8277 (
            .O(N__38521),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__8276 (
            .O(N__38518),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8275 (
            .O(N__38513),
            .I(N__38510));
    LocalMux I__8274 (
            .O(N__38510),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    InMux I__8273 (
            .O(N__38507),
            .I(N__38503));
    InMux I__8272 (
            .O(N__38506),
            .I(N__38500));
    LocalMux I__8271 (
            .O(N__38503),
            .I(N__38497));
    LocalMux I__8270 (
            .O(N__38500),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__8269 (
            .O(N__38497),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8268 (
            .O(N__38492),
            .I(N__38489));
    LocalMux I__8267 (
            .O(N__38489),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    InMux I__8266 (
            .O(N__38486),
            .I(N__38482));
    InMux I__8265 (
            .O(N__38485),
            .I(N__38479));
    LocalMux I__8264 (
            .O(N__38482),
            .I(N__38476));
    LocalMux I__8263 (
            .O(N__38479),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__8262 (
            .O(N__38476),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8261 (
            .O(N__38471),
            .I(N__38468));
    LocalMux I__8260 (
            .O(N__38468),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    InMux I__8259 (
            .O(N__38465),
            .I(N__38461));
    InMux I__8258 (
            .O(N__38464),
            .I(N__38458));
    LocalMux I__8257 (
            .O(N__38461),
            .I(N__38455));
    LocalMux I__8256 (
            .O(N__38458),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__8255 (
            .O(N__38455),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8254 (
            .O(N__38450),
            .I(N__38447));
    LocalMux I__8253 (
            .O(N__38447),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    InMux I__8252 (
            .O(N__38444),
            .I(N__38440));
    InMux I__8251 (
            .O(N__38443),
            .I(N__38437));
    LocalMux I__8250 (
            .O(N__38440),
            .I(N__38434));
    LocalMux I__8249 (
            .O(N__38437),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__8248 (
            .O(N__38434),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__8247 (
            .O(N__38429),
            .I(N__38426));
    InMux I__8246 (
            .O(N__38426),
            .I(N__38423));
    LocalMux I__8245 (
            .O(N__38423),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__8244 (
            .O(N__38420),
            .I(N__38417));
    InMux I__8243 (
            .O(N__38417),
            .I(N__38414));
    LocalMux I__8242 (
            .O(N__38414),
            .I(N__38411));
    Odrv12 I__8241 (
            .O(N__38411),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    InMux I__8240 (
            .O(N__38408),
            .I(N__38404));
    CascadeMux I__8239 (
            .O(N__38407),
            .I(N__38401));
    LocalMux I__8238 (
            .O(N__38404),
            .I(N__38398));
    InMux I__8237 (
            .O(N__38401),
            .I(N__38395));
    Span4Mux_v I__8236 (
            .O(N__38398),
            .I(N__38392));
    LocalMux I__8235 (
            .O(N__38395),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8234 (
            .O(N__38392),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__8233 (
            .O(N__38387),
            .I(N__38384));
    LocalMux I__8232 (
            .O(N__38384),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    InMux I__8231 (
            .O(N__38381),
            .I(N__38378));
    LocalMux I__8230 (
            .O(N__38378),
            .I(N__38374));
    InMux I__8229 (
            .O(N__38377),
            .I(N__38371));
    Odrv4 I__8228 (
            .O(N__38374),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__8227 (
            .O(N__38371),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8226 (
            .O(N__38366),
            .I(N__38363));
    LocalMux I__8225 (
            .O(N__38363),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__8224 (
            .O(N__38360),
            .I(N__38357));
    InMux I__8223 (
            .O(N__38357),
            .I(N__38354));
    LocalMux I__8222 (
            .O(N__38354),
            .I(N__38350));
    InMux I__8221 (
            .O(N__38353),
            .I(N__38347));
    Odrv4 I__8220 (
            .O(N__38350),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__8219 (
            .O(N__38347),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8218 (
            .O(N__38342),
            .I(N__38339));
    LocalMux I__8217 (
            .O(N__38339),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    InMux I__8216 (
            .O(N__38336),
            .I(N__38333));
    LocalMux I__8215 (
            .O(N__38333),
            .I(N__38329));
    InMux I__8214 (
            .O(N__38332),
            .I(N__38326));
    Odrv4 I__8213 (
            .O(N__38329),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__8212 (
            .O(N__38326),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8211 (
            .O(N__38321),
            .I(N__38318));
    LocalMux I__8210 (
            .O(N__38318),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    InMux I__8209 (
            .O(N__38315),
            .I(N__38312));
    LocalMux I__8208 (
            .O(N__38312),
            .I(N__38308));
    InMux I__8207 (
            .O(N__38311),
            .I(N__38305));
    Odrv12 I__8206 (
            .O(N__38308),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__8205 (
            .O(N__38305),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8204 (
            .O(N__38300),
            .I(N__38297));
    LocalMux I__8203 (
            .O(N__38297),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__8202 (
            .O(N__38294),
            .I(N__38291));
    InMux I__8201 (
            .O(N__38291),
            .I(N__38288));
    LocalMux I__8200 (
            .O(N__38288),
            .I(N__38284));
    InMux I__8199 (
            .O(N__38287),
            .I(N__38281));
    Odrv12 I__8198 (
            .O(N__38284),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__8197 (
            .O(N__38281),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8196 (
            .O(N__38276),
            .I(N__38273));
    LocalMux I__8195 (
            .O(N__38273),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    InMux I__8194 (
            .O(N__38270),
            .I(N__38266));
    InMux I__8193 (
            .O(N__38269),
            .I(N__38263));
    LocalMux I__8192 (
            .O(N__38266),
            .I(N__38260));
    LocalMux I__8191 (
            .O(N__38263),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__8190 (
            .O(N__38260),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8189 (
            .O(N__38255),
            .I(N__38252));
    LocalMux I__8188 (
            .O(N__38252),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__8187 (
            .O(N__38249),
            .I(N__38246));
    InMux I__8186 (
            .O(N__38246),
            .I(N__38243));
    LocalMux I__8185 (
            .O(N__38243),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    InMux I__8184 (
            .O(N__38240),
            .I(N__38236));
    InMux I__8183 (
            .O(N__38239),
            .I(N__38233));
    LocalMux I__8182 (
            .O(N__38236),
            .I(N__38230));
    LocalMux I__8181 (
            .O(N__38233),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__8180 (
            .O(N__38230),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8179 (
            .O(N__38225),
            .I(N__38222));
    LocalMux I__8178 (
            .O(N__38222),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    InMux I__8177 (
            .O(N__38219),
            .I(N__38215));
    InMux I__8176 (
            .O(N__38218),
            .I(N__38212));
    LocalMux I__8175 (
            .O(N__38215),
            .I(N__38209));
    LocalMux I__8174 (
            .O(N__38212),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__8173 (
            .O(N__38209),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8172 (
            .O(N__38204),
            .I(N__38201));
    LocalMux I__8171 (
            .O(N__38201),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    InMux I__8170 (
            .O(N__38198),
            .I(N__38195));
    LocalMux I__8169 (
            .O(N__38195),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__8168 (
            .O(N__38192),
            .I(N__38186));
    InMux I__8167 (
            .O(N__38191),
            .I(N__38183));
    InMux I__8166 (
            .O(N__38190),
            .I(N__38180));
    InMux I__8165 (
            .O(N__38189),
            .I(N__38177));
    LocalMux I__8164 (
            .O(N__38186),
            .I(N__38170));
    LocalMux I__8163 (
            .O(N__38183),
            .I(N__38170));
    LocalMux I__8162 (
            .O(N__38180),
            .I(N__38170));
    LocalMux I__8161 (
            .O(N__38177),
            .I(N__38167));
    Span4Mux_v I__8160 (
            .O(N__38170),
            .I(N__38164));
    Odrv4 I__8159 (
            .O(N__38167),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    Odrv4 I__8158 (
            .O(N__38164),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    CascadeMux I__8157 (
            .O(N__38159),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__8156 (
            .O(N__38156),
            .I(N__38153));
    LocalMux I__8155 (
            .O(N__38153),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__8154 (
            .O(N__38150),
            .I(N__38147));
    LocalMux I__8153 (
            .O(N__38147),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__8152 (
            .O(N__38144),
            .I(N__38141));
    LocalMux I__8151 (
            .O(N__38141),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__8150 (
            .O(N__38138),
            .I(N__38135));
    LocalMux I__8149 (
            .O(N__38135),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    CascadeMux I__8148 (
            .O(N__38132),
            .I(N__38126));
    CascadeMux I__8147 (
            .O(N__38131),
            .I(N__38110));
    CascadeMux I__8146 (
            .O(N__38130),
            .I(N__38107));
    InMux I__8145 (
            .O(N__38129),
            .I(N__38089));
    InMux I__8144 (
            .O(N__38126),
            .I(N__38089));
    InMux I__8143 (
            .O(N__38125),
            .I(N__38089));
    InMux I__8142 (
            .O(N__38124),
            .I(N__38089));
    InMux I__8141 (
            .O(N__38123),
            .I(N__38089));
    InMux I__8140 (
            .O(N__38122),
            .I(N__38089));
    InMux I__8139 (
            .O(N__38121),
            .I(N__38089));
    InMux I__8138 (
            .O(N__38120),
            .I(N__38072));
    InMux I__8137 (
            .O(N__38119),
            .I(N__38072));
    InMux I__8136 (
            .O(N__38118),
            .I(N__38072));
    InMux I__8135 (
            .O(N__38117),
            .I(N__38072));
    InMux I__8134 (
            .O(N__38116),
            .I(N__38072));
    InMux I__8133 (
            .O(N__38115),
            .I(N__38072));
    InMux I__8132 (
            .O(N__38114),
            .I(N__38072));
    InMux I__8131 (
            .O(N__38113),
            .I(N__38072));
    InMux I__8130 (
            .O(N__38110),
            .I(N__38063));
    InMux I__8129 (
            .O(N__38107),
            .I(N__38063));
    InMux I__8128 (
            .O(N__38106),
            .I(N__38063));
    InMux I__8127 (
            .O(N__38105),
            .I(N__38063));
    CascadeMux I__8126 (
            .O(N__38104),
            .I(N__38059));
    LocalMux I__8125 (
            .O(N__38089),
            .I(N__38055));
    LocalMux I__8124 (
            .O(N__38072),
            .I(N__38052));
    LocalMux I__8123 (
            .O(N__38063),
            .I(N__38049));
    InMux I__8122 (
            .O(N__38062),
            .I(N__38042));
    InMux I__8121 (
            .O(N__38059),
            .I(N__38042));
    InMux I__8120 (
            .O(N__38058),
            .I(N__38039));
    Span4Mux_v I__8119 (
            .O(N__38055),
            .I(N__38034));
    Span4Mux_v I__8118 (
            .O(N__38052),
            .I(N__38034));
    Span4Mux_h I__8117 (
            .O(N__38049),
            .I(N__38031));
    InMux I__8116 (
            .O(N__38048),
            .I(N__38026));
    InMux I__8115 (
            .O(N__38047),
            .I(N__38026));
    LocalMux I__8114 (
            .O(N__38042),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__8113 (
            .O(N__38039),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__8112 (
            .O(N__38034),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__8111 (
            .O(N__38031),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__8110 (
            .O(N__38026),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__8109 (
            .O(N__38015),
            .I(N__38004));
    CascadeMux I__8108 (
            .O(N__38014),
            .I(N__38001));
    CascadeMux I__8107 (
            .O(N__38013),
            .I(N__37998));
    CascadeMux I__8106 (
            .O(N__38012),
            .I(N__37995));
    CascadeMux I__8105 (
            .O(N__38011),
            .I(N__37988));
    CascadeMux I__8104 (
            .O(N__38010),
            .I(N__37985));
    CascadeMux I__8103 (
            .O(N__38009),
            .I(N__37982));
    CascadeMux I__8102 (
            .O(N__38008),
            .I(N__37975));
    InMux I__8101 (
            .O(N__38007),
            .I(N__37969));
    InMux I__8100 (
            .O(N__38004),
            .I(N__37952));
    InMux I__8099 (
            .O(N__38001),
            .I(N__37952));
    InMux I__8098 (
            .O(N__37998),
            .I(N__37952));
    InMux I__8097 (
            .O(N__37995),
            .I(N__37952));
    InMux I__8096 (
            .O(N__37994),
            .I(N__37952));
    InMux I__8095 (
            .O(N__37993),
            .I(N__37952));
    InMux I__8094 (
            .O(N__37992),
            .I(N__37952));
    InMux I__8093 (
            .O(N__37991),
            .I(N__37952));
    InMux I__8092 (
            .O(N__37988),
            .I(N__37939));
    InMux I__8091 (
            .O(N__37985),
            .I(N__37939));
    InMux I__8090 (
            .O(N__37982),
            .I(N__37939));
    InMux I__8089 (
            .O(N__37981),
            .I(N__37939));
    InMux I__8088 (
            .O(N__37980),
            .I(N__37939));
    InMux I__8087 (
            .O(N__37979),
            .I(N__37939));
    CascadeMux I__8086 (
            .O(N__37978),
            .I(N__37935));
    InMux I__8085 (
            .O(N__37975),
            .I(N__37928));
    InMux I__8084 (
            .O(N__37974),
            .I(N__37928));
    InMux I__8083 (
            .O(N__37973),
            .I(N__37925));
    CascadeMux I__8082 (
            .O(N__37972),
            .I(N__37922));
    LocalMux I__8081 (
            .O(N__37969),
            .I(N__37914));
    LocalMux I__8080 (
            .O(N__37952),
            .I(N__37914));
    LocalMux I__8079 (
            .O(N__37939),
            .I(N__37914));
    InMux I__8078 (
            .O(N__37938),
            .I(N__37905));
    InMux I__8077 (
            .O(N__37935),
            .I(N__37905));
    InMux I__8076 (
            .O(N__37934),
            .I(N__37905));
    InMux I__8075 (
            .O(N__37933),
            .I(N__37905));
    LocalMux I__8074 (
            .O(N__37928),
            .I(N__37900));
    LocalMux I__8073 (
            .O(N__37925),
            .I(N__37900));
    InMux I__8072 (
            .O(N__37922),
            .I(N__37897));
    InMux I__8071 (
            .O(N__37921),
            .I(N__37894));
    Span4Mux_v I__8070 (
            .O(N__37914),
            .I(N__37891));
    LocalMux I__8069 (
            .O(N__37905),
            .I(N__37888));
    Span4Mux_v I__8068 (
            .O(N__37900),
            .I(N__37885));
    LocalMux I__8067 (
            .O(N__37897),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__8066 (
            .O(N__37894),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__8065 (
            .O(N__37891),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__8064 (
            .O(N__37888),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__8063 (
            .O(N__37885),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    CascadeMux I__8062 (
            .O(N__37874),
            .I(N__37866));
    CascadeMux I__8061 (
            .O(N__37873),
            .I(N__37863));
    CascadeMux I__8060 (
            .O(N__37872),
            .I(N__37855));
    CascadeMux I__8059 (
            .O(N__37871),
            .I(N__37852));
    CascadeMux I__8058 (
            .O(N__37870),
            .I(N__37849));
    CascadeMux I__8057 (
            .O(N__37869),
            .I(N__37846));
    InMux I__8056 (
            .O(N__37866),
            .I(N__37833));
    InMux I__8055 (
            .O(N__37863),
            .I(N__37833));
    InMux I__8054 (
            .O(N__37862),
            .I(N__37822));
    InMux I__8053 (
            .O(N__37861),
            .I(N__37822));
    InMux I__8052 (
            .O(N__37860),
            .I(N__37822));
    InMux I__8051 (
            .O(N__37859),
            .I(N__37822));
    InMux I__8050 (
            .O(N__37858),
            .I(N__37822));
    InMux I__8049 (
            .O(N__37855),
            .I(N__37813));
    InMux I__8048 (
            .O(N__37852),
            .I(N__37813));
    InMux I__8047 (
            .O(N__37849),
            .I(N__37813));
    InMux I__8046 (
            .O(N__37846),
            .I(N__37813));
    InMux I__8045 (
            .O(N__37845),
            .I(N__37804));
    InMux I__8044 (
            .O(N__37844),
            .I(N__37804));
    InMux I__8043 (
            .O(N__37843),
            .I(N__37804));
    InMux I__8042 (
            .O(N__37842),
            .I(N__37804));
    InMux I__8041 (
            .O(N__37841),
            .I(N__37799));
    InMux I__8040 (
            .O(N__37840),
            .I(N__37799));
    InMux I__8039 (
            .O(N__37839),
            .I(N__37794));
    InMux I__8038 (
            .O(N__37838),
            .I(N__37794));
    LocalMux I__8037 (
            .O(N__37833),
            .I(N__37786));
    LocalMux I__8036 (
            .O(N__37822),
            .I(N__37786));
    LocalMux I__8035 (
            .O(N__37813),
            .I(N__37781));
    LocalMux I__8034 (
            .O(N__37804),
            .I(N__37781));
    LocalMux I__8033 (
            .O(N__37799),
            .I(N__37775));
    LocalMux I__8032 (
            .O(N__37794),
            .I(N__37775));
    InMux I__8031 (
            .O(N__37793),
            .I(N__37769));
    InMux I__8030 (
            .O(N__37792),
            .I(N__37769));
    InMux I__8029 (
            .O(N__37791),
            .I(N__37766));
    Span4Mux_h I__8028 (
            .O(N__37786),
            .I(N__37761));
    Span4Mux_v I__8027 (
            .O(N__37781),
            .I(N__37761));
    InMux I__8026 (
            .O(N__37780),
            .I(N__37758));
    Span4Mux_h I__8025 (
            .O(N__37775),
            .I(N__37755));
    InMux I__8024 (
            .O(N__37774),
            .I(N__37752));
    LocalMux I__8023 (
            .O(N__37769),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__8022 (
            .O(N__37766),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__8021 (
            .O(N__37761),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__8020 (
            .O(N__37758),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__8019 (
            .O(N__37755),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__8018 (
            .O(N__37752),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__8017 (
            .O(N__37739),
            .I(N__37736));
    LocalMux I__8016 (
            .O(N__37736),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    CascadeMux I__8015 (
            .O(N__37733),
            .I(N__37730));
    InMux I__8014 (
            .O(N__37730),
            .I(N__37726));
    InMux I__8013 (
            .O(N__37729),
            .I(N__37722));
    LocalMux I__8012 (
            .O(N__37726),
            .I(N__37719));
    InMux I__8011 (
            .O(N__37725),
            .I(N__37716));
    LocalMux I__8010 (
            .O(N__37722),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__8009 (
            .O(N__37719),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8008 (
            .O(N__37716),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8007 (
            .O(N__37709),
            .I(N__37706));
    LocalMux I__8006 (
            .O(N__37706),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    InMux I__8005 (
            .O(N__37703),
            .I(N__37700));
    LocalMux I__8004 (
            .O(N__37700),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__8003 (
            .O(N__37697),
            .I(N__37694));
    InMux I__8002 (
            .O(N__37694),
            .I(N__37691));
    LocalMux I__8001 (
            .O(N__37691),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__8000 (
            .O(N__37688),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__7999 (
            .O(N__37685),
            .I(N__37682));
    LocalMux I__7998 (
            .O(N__37682),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ));
    InMux I__7997 (
            .O(N__37679),
            .I(N__37676));
    LocalMux I__7996 (
            .O(N__37676),
            .I(N__37673));
    Span4Mux_v I__7995 (
            .O(N__37673),
            .I(N__37670));
    Odrv4 I__7994 (
            .O(N__37670),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    InMux I__7993 (
            .O(N__37667),
            .I(N__37664));
    LocalMux I__7992 (
            .O(N__37664),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__7991 (
            .O(N__37661),
            .I(N__37658));
    LocalMux I__7990 (
            .O(N__37658),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__7989 (
            .O(N__37655),
            .I(N__37652));
    LocalMux I__7988 (
            .O(N__37652),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__7987 (
            .O(N__37649),
            .I(N__37646));
    LocalMux I__7986 (
            .O(N__37646),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    CascadeMux I__7985 (
            .O(N__37643),
            .I(N__37640));
    InMux I__7984 (
            .O(N__37640),
            .I(N__37637));
    LocalMux I__7983 (
            .O(N__37637),
            .I(N__37634));
    Span4Mux_h I__7982 (
            .O(N__37634),
            .I(N__37631));
    Odrv4 I__7981 (
            .O(N__37631),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    InMux I__7980 (
            .O(N__37628),
            .I(N__37625));
    LocalMux I__7979 (
            .O(N__37625),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__7978 (
            .O(N__37622),
            .I(N__37619));
    InMux I__7977 (
            .O(N__37619),
            .I(N__37616));
    LocalMux I__7976 (
            .O(N__37616),
            .I(N__37613));
    Odrv4 I__7975 (
            .O(N__37613),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__7974 (
            .O(N__37610),
            .I(N__37607));
    LocalMux I__7973 (
            .O(N__37607),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__7972 (
            .O(N__37604),
            .I(N__37601));
    InMux I__7971 (
            .O(N__37601),
            .I(N__37598));
    LocalMux I__7970 (
            .O(N__37598),
            .I(N__37595));
    Odrv4 I__7969 (
            .O(N__37595),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    InMux I__7968 (
            .O(N__37592),
            .I(N__37589));
    LocalMux I__7967 (
            .O(N__37589),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__7966 (
            .O(N__37586),
            .I(N__37583));
    InMux I__7965 (
            .O(N__37583),
            .I(N__37580));
    LocalMux I__7964 (
            .O(N__37580),
            .I(N__37577));
    Span4Mux_v I__7963 (
            .O(N__37577),
            .I(N__37574));
    Odrv4 I__7962 (
            .O(N__37574),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__7961 (
            .O(N__37571),
            .I(N__37568));
    LocalMux I__7960 (
            .O(N__37568),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__7959 (
            .O(N__37565),
            .I(N__37562));
    InMux I__7958 (
            .O(N__37562),
            .I(N__37559));
    LocalMux I__7957 (
            .O(N__37559),
            .I(N__37556));
    Odrv4 I__7956 (
            .O(N__37556),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__7955 (
            .O(N__37553),
            .I(N__37550));
    LocalMux I__7954 (
            .O(N__37550),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__7953 (
            .O(N__37547),
            .I(N__37544));
    InMux I__7952 (
            .O(N__37544),
            .I(N__37541));
    LocalMux I__7951 (
            .O(N__37541),
            .I(N__37538));
    Span4Mux_h I__7950 (
            .O(N__37538),
            .I(N__37535));
    Odrv4 I__7949 (
            .O(N__37535),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__7948 (
            .O(N__37532),
            .I(N__37529));
    LocalMux I__7947 (
            .O(N__37529),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__7946 (
            .O(N__37526),
            .I(N__37523));
    InMux I__7945 (
            .O(N__37523),
            .I(N__37520));
    LocalMux I__7944 (
            .O(N__37520),
            .I(N__37517));
    Span4Mux_h I__7943 (
            .O(N__37517),
            .I(N__37514));
    Odrv4 I__7942 (
            .O(N__37514),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    InMux I__7941 (
            .O(N__37511),
            .I(N__37508));
    LocalMux I__7940 (
            .O(N__37508),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__7939 (
            .O(N__37505),
            .I(N__37502));
    InMux I__7938 (
            .O(N__37502),
            .I(N__37499));
    LocalMux I__7937 (
            .O(N__37499),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    InMux I__7936 (
            .O(N__37496),
            .I(N__37493));
    LocalMux I__7935 (
            .O(N__37493),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__7934 (
            .O(N__37490),
            .I(N__37487));
    InMux I__7933 (
            .O(N__37487),
            .I(N__37484));
    LocalMux I__7932 (
            .O(N__37484),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__7931 (
            .O(N__37481),
            .I(N__37478));
    LocalMux I__7930 (
            .O(N__37478),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__7929 (
            .O(N__37475),
            .I(N__37472));
    InMux I__7928 (
            .O(N__37472),
            .I(N__37469));
    LocalMux I__7927 (
            .O(N__37469),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    InMux I__7926 (
            .O(N__37466),
            .I(N__37463));
    LocalMux I__7925 (
            .O(N__37463),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__7924 (
            .O(N__37460),
            .I(N__37457));
    InMux I__7923 (
            .O(N__37457),
            .I(N__37454));
    LocalMux I__7922 (
            .O(N__37454),
            .I(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ));
    InMux I__7921 (
            .O(N__37451),
            .I(N__37448));
    LocalMux I__7920 (
            .O(N__37448),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__7919 (
            .O(N__37445),
            .I(N__37442));
    InMux I__7918 (
            .O(N__37442),
            .I(N__37439));
    LocalMux I__7917 (
            .O(N__37439),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__7916 (
            .O(N__37436),
            .I(N__37433));
    LocalMux I__7915 (
            .O(N__37433),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__7914 (
            .O(N__37430),
            .I(N__37427));
    InMux I__7913 (
            .O(N__37427),
            .I(N__37424));
    LocalMux I__7912 (
            .O(N__37424),
            .I(N__37421));
    Odrv12 I__7911 (
            .O(N__37421),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    InMux I__7910 (
            .O(N__37418),
            .I(N__37415));
    LocalMux I__7909 (
            .O(N__37415),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__7908 (
            .O(N__37412),
            .I(N__37409));
    InMux I__7907 (
            .O(N__37409),
            .I(N__37406));
    LocalMux I__7906 (
            .O(N__37406),
            .I(N__37403));
    Odrv4 I__7905 (
            .O(N__37403),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    InMux I__7904 (
            .O(N__37400),
            .I(N__37397));
    LocalMux I__7903 (
            .O(N__37397),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__7902 (
            .O(N__37394),
            .I(N__37391));
    InMux I__7901 (
            .O(N__37391),
            .I(N__37388));
    LocalMux I__7900 (
            .O(N__37388),
            .I(N__37385));
    Odrv4 I__7899 (
            .O(N__37385),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__7898 (
            .O(N__37382),
            .I(N__37379));
    LocalMux I__7897 (
            .O(N__37379),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    InMux I__7896 (
            .O(N__37376),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__7895 (
            .O(N__37373),
            .I(N__37369));
    InMux I__7894 (
            .O(N__37372),
            .I(N__37366));
    LocalMux I__7893 (
            .O(N__37369),
            .I(N__37363));
    LocalMux I__7892 (
            .O(N__37366),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__7891 (
            .O(N__37363),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__7890 (
            .O(N__37358),
            .I(N__37355));
    InMux I__7889 (
            .O(N__37355),
            .I(N__37352));
    LocalMux I__7888 (
            .O(N__37352),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__7887 (
            .O(N__37349),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__7886 (
            .O(N__37346),
            .I(N__37342));
    InMux I__7885 (
            .O(N__37345),
            .I(N__37339));
    LocalMux I__7884 (
            .O(N__37342),
            .I(N__37336));
    LocalMux I__7883 (
            .O(N__37339),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__7882 (
            .O(N__37336),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__7881 (
            .O(N__37331),
            .I(N__37328));
    LocalMux I__7880 (
            .O(N__37328),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__7879 (
            .O(N__37325),
            .I(bfn_15_15_0_));
    InMux I__7878 (
            .O(N__37322),
            .I(N__37318));
    InMux I__7877 (
            .O(N__37321),
            .I(N__37315));
    LocalMux I__7876 (
            .O(N__37318),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__7875 (
            .O(N__37315),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__7874 (
            .O(N__37310),
            .I(N__37307));
    InMux I__7873 (
            .O(N__37307),
            .I(N__37304));
    LocalMux I__7872 (
            .O(N__37304),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__7871 (
            .O(N__37301),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__7870 (
            .O(N__37298),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    CascadeMux I__7869 (
            .O(N__37295),
            .I(N__37292));
    InMux I__7868 (
            .O(N__37292),
            .I(N__37289));
    LocalMux I__7867 (
            .O(N__37289),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__7866 (
            .O(N__37286),
            .I(N__37283));
    InMux I__7865 (
            .O(N__37283),
            .I(N__37280));
    LocalMux I__7864 (
            .O(N__37280),
            .I(N__37277));
    Odrv4 I__7863 (
            .O(N__37277),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    InMux I__7862 (
            .O(N__37274),
            .I(N__37271));
    LocalMux I__7861 (
            .O(N__37271),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__7860 (
            .O(N__37268),
            .I(N__37265));
    InMux I__7859 (
            .O(N__37265),
            .I(N__37262));
    LocalMux I__7858 (
            .O(N__37262),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__7857 (
            .O(N__37259),
            .I(N__37256));
    LocalMux I__7856 (
            .O(N__37256),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__7855 (
            .O(N__37253),
            .I(N__37250));
    InMux I__7854 (
            .O(N__37250),
            .I(N__37247));
    LocalMux I__7853 (
            .O(N__37247),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    InMux I__7852 (
            .O(N__37244),
            .I(N__37241));
    LocalMux I__7851 (
            .O(N__37241),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    InMux I__7850 (
            .O(N__37238),
            .I(N__37235));
    LocalMux I__7849 (
            .O(N__37235),
            .I(N__37232));
    Span4Mux_h I__7848 (
            .O(N__37232),
            .I(N__37228));
    InMux I__7847 (
            .O(N__37231),
            .I(N__37225));
    Odrv4 I__7846 (
            .O(N__37228),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__7845 (
            .O(N__37225),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__7844 (
            .O(N__37220),
            .I(N__37217));
    LocalMux I__7843 (
            .O(N__37217),
            .I(N__37214));
    Span4Mux_h I__7842 (
            .O(N__37214),
            .I(N__37211));
    Odrv4 I__7841 (
            .O(N__37211),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__7840 (
            .O(N__37208),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__7839 (
            .O(N__37205),
            .I(N__37201));
    InMux I__7838 (
            .O(N__37204),
            .I(N__37198));
    LocalMux I__7837 (
            .O(N__37201),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__7836 (
            .O(N__37198),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__7835 (
            .O(N__37193),
            .I(N__37190));
    InMux I__7834 (
            .O(N__37190),
            .I(N__37187));
    LocalMux I__7833 (
            .O(N__37187),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__7832 (
            .O(N__37184),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__7831 (
            .O(N__37181),
            .I(N__37178));
    LocalMux I__7830 (
            .O(N__37178),
            .I(N__37174));
    InMux I__7829 (
            .O(N__37177),
            .I(N__37171));
    Odrv4 I__7828 (
            .O(N__37174),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__7827 (
            .O(N__37171),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__7826 (
            .O(N__37166),
            .I(N__37163));
    LocalMux I__7825 (
            .O(N__37163),
            .I(N__37160));
    Odrv12 I__7824 (
            .O(N__37160),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__7823 (
            .O(N__37157),
            .I(bfn_15_14_0_));
    InMux I__7822 (
            .O(N__37154),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__7821 (
            .O(N__37151),
            .I(N__37148));
    LocalMux I__7820 (
            .O(N__37148),
            .I(N__37144));
    InMux I__7819 (
            .O(N__37147),
            .I(N__37141));
    Odrv4 I__7818 (
            .O(N__37144),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__7817 (
            .O(N__37141),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__7816 (
            .O(N__37136),
            .I(N__37133));
    InMux I__7815 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7814 (
            .O(N__37130),
            .I(N__37127));
    Odrv4 I__7813 (
            .O(N__37127),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__7812 (
            .O(N__37124),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__7811 (
            .O(N__37121),
            .I(N__37117));
    InMux I__7810 (
            .O(N__37120),
            .I(N__37114));
    LocalMux I__7809 (
            .O(N__37117),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__7808 (
            .O(N__37114),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__7807 (
            .O(N__37109),
            .I(N__37106));
    LocalMux I__7806 (
            .O(N__37106),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__7805 (
            .O(N__37103),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__7804 (
            .O(N__37100),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__7803 (
            .O(N__37097),
            .I(N__37093));
    InMux I__7802 (
            .O(N__37096),
            .I(N__37090));
    LocalMux I__7801 (
            .O(N__37093),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__7800 (
            .O(N__37090),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__7799 (
            .O(N__37085),
            .I(N__37082));
    LocalMux I__7798 (
            .O(N__37082),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__7797 (
            .O(N__37079),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__7796 (
            .O(N__37076),
            .I(N__37072));
    InMux I__7795 (
            .O(N__37075),
            .I(N__37069));
    LocalMux I__7794 (
            .O(N__37072),
            .I(measured_delay_hc_29));
    LocalMux I__7793 (
            .O(N__37069),
            .I(measured_delay_hc_29));
    InMux I__7792 (
            .O(N__37064),
            .I(N__37061));
    LocalMux I__7791 (
            .O(N__37061),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ));
    CascadeMux I__7790 (
            .O(N__37058),
            .I(N__37054));
    InMux I__7789 (
            .O(N__37057),
            .I(N__37051));
    InMux I__7788 (
            .O(N__37054),
            .I(N__37048));
    LocalMux I__7787 (
            .O(N__37051),
            .I(measured_delay_hc_27));
    LocalMux I__7786 (
            .O(N__37048),
            .I(measured_delay_hc_27));
    InMux I__7785 (
            .O(N__37043),
            .I(N__37040));
    LocalMux I__7784 (
            .O(N__37040),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    CascadeMux I__7783 (
            .O(N__37037),
            .I(N__37034));
    InMux I__7782 (
            .O(N__37034),
            .I(N__37031));
    LocalMux I__7781 (
            .O(N__37031),
            .I(N__37027));
    InMux I__7780 (
            .O(N__37030),
            .I(N__37023));
    Span4Mux_h I__7779 (
            .O(N__37027),
            .I(N__37020));
    InMux I__7778 (
            .O(N__37026),
            .I(N__37017));
    LocalMux I__7777 (
            .O(N__37023),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7776 (
            .O(N__37020),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__7775 (
            .O(N__37017),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__7774 (
            .O(N__37010),
            .I(N__37006));
    InMux I__7773 (
            .O(N__37009),
            .I(N__37003));
    LocalMux I__7772 (
            .O(N__37006),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__7771 (
            .O(N__37003),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__7770 (
            .O(N__36998),
            .I(N__36995));
    InMux I__7769 (
            .O(N__36995),
            .I(N__36992));
    LocalMux I__7768 (
            .O(N__36992),
            .I(N__36989));
    Span4Mux_h I__7767 (
            .O(N__36989),
            .I(N__36986));
    Odrv4 I__7766 (
            .O(N__36986),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__7765 (
            .O(N__36983),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__7764 (
            .O(N__36980),
            .I(N__36977));
    LocalMux I__7763 (
            .O(N__36977),
            .I(N__36974));
    Span4Mux_v I__7762 (
            .O(N__36974),
            .I(N__36971));
    Odrv4 I__7761 (
            .O(N__36971),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    CascadeMux I__7760 (
            .O(N__36968),
            .I(N__36965));
    InMux I__7759 (
            .O(N__36965),
            .I(N__36961));
    InMux I__7758 (
            .O(N__36964),
            .I(N__36958));
    LocalMux I__7757 (
            .O(N__36961),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__7756 (
            .O(N__36958),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__7755 (
            .O(N__36953),
            .I(N__36950));
    LocalMux I__7754 (
            .O(N__36950),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__7753 (
            .O(N__36947),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__7752 (
            .O(N__36944),
            .I(N__36941));
    LocalMux I__7751 (
            .O(N__36941),
            .I(N__36938));
    Span4Mux_v I__7750 (
            .O(N__36938),
            .I(N__36934));
    InMux I__7749 (
            .O(N__36937),
            .I(N__36931));
    Odrv4 I__7748 (
            .O(N__36934),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__7747 (
            .O(N__36931),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__7746 (
            .O(N__36926),
            .I(N__36923));
    InMux I__7745 (
            .O(N__36923),
            .I(N__36920));
    LocalMux I__7744 (
            .O(N__36920),
            .I(N__36917));
    Span4Mux_h I__7743 (
            .O(N__36917),
            .I(N__36914));
    Odrv4 I__7742 (
            .O(N__36914),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__7741 (
            .O(N__36911),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__7740 (
            .O(N__36908),
            .I(N__36905));
    LocalMux I__7739 (
            .O(N__36905),
            .I(N__36902));
    Span4Mux_h I__7738 (
            .O(N__36902),
            .I(N__36898));
    InMux I__7737 (
            .O(N__36901),
            .I(N__36895));
    Odrv4 I__7736 (
            .O(N__36898),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__7735 (
            .O(N__36895),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__7734 (
            .O(N__36890),
            .I(N__36887));
    LocalMux I__7733 (
            .O(N__36887),
            .I(N__36884));
    Span4Mux_v I__7732 (
            .O(N__36884),
            .I(N__36881));
    Odrv4 I__7731 (
            .O(N__36881),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__7730 (
            .O(N__36878),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__7729 (
            .O(N__36875),
            .I(N__36871));
    InMux I__7728 (
            .O(N__36874),
            .I(N__36868));
    LocalMux I__7727 (
            .O(N__36871),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__7726 (
            .O(N__36868),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__7725 (
            .O(N__36863),
            .I(N__36860));
    InMux I__7724 (
            .O(N__36860),
            .I(N__36857));
    LocalMux I__7723 (
            .O(N__36857),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__7722 (
            .O(N__36854),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    CascadeMux I__7721 (
            .O(N__36851),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_c_cascade_ ));
    CascadeMux I__7720 (
            .O(N__36848),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_0_0_cascade_ ));
    InMux I__7719 (
            .O(N__36845),
            .I(N__36842));
    LocalMux I__7718 (
            .O(N__36842),
            .I(N__36839));
    Span12Mux_v I__7717 (
            .O(N__36839),
            .I(N__36836));
    Odrv12 I__7716 (
            .O(N__36836),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13 ));
    CascadeMux I__7715 (
            .O(N__36833),
            .I(N__36830));
    InMux I__7714 (
            .O(N__36830),
            .I(N__36827));
    LocalMux I__7713 (
            .O(N__36827),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9 ));
    InMux I__7712 (
            .O(N__36824),
            .I(N__36820));
    InMux I__7711 (
            .O(N__36823),
            .I(N__36816));
    LocalMux I__7710 (
            .O(N__36820),
            .I(N__36813));
    InMux I__7709 (
            .O(N__36819),
            .I(N__36810));
    LocalMux I__7708 (
            .O(N__36816),
            .I(N__36805));
    Span12Mux_s10_h I__7707 (
            .O(N__36813),
            .I(N__36805));
    LocalMux I__7706 (
            .O(N__36810),
            .I(measured_delay_hc_21));
    Odrv12 I__7705 (
            .O(N__36805),
            .I(measured_delay_hc_21));
    InMux I__7704 (
            .O(N__36800),
            .I(N__36796));
    InMux I__7703 (
            .O(N__36799),
            .I(N__36793));
    LocalMux I__7702 (
            .O(N__36796),
            .I(N__36789));
    LocalMux I__7701 (
            .O(N__36793),
            .I(N__36786));
    InMux I__7700 (
            .O(N__36792),
            .I(N__36783));
    Span12Mux_v I__7699 (
            .O(N__36789),
            .I(N__36780));
    Span4Mux_v I__7698 (
            .O(N__36786),
            .I(N__36777));
    LocalMux I__7697 (
            .O(N__36783),
            .I(N__36774));
    Odrv12 I__7696 (
            .O(N__36780),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    Odrv4 I__7695 (
            .O(N__36777),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    Odrv4 I__7694 (
            .O(N__36774),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    CascadeMux I__7693 (
            .O(N__36767),
            .I(N__36764));
    InMux I__7692 (
            .O(N__36764),
            .I(N__36759));
    InMux I__7691 (
            .O(N__36763),
            .I(N__36754));
    InMux I__7690 (
            .O(N__36762),
            .I(N__36754));
    LocalMux I__7689 (
            .O(N__36759),
            .I(N__36751));
    LocalMux I__7688 (
            .O(N__36754),
            .I(measured_delay_hc_20));
    Odrv4 I__7687 (
            .O(N__36751),
            .I(measured_delay_hc_20));
    CascadeMux I__7686 (
            .O(N__36746),
            .I(N__36743));
    InMux I__7685 (
            .O(N__36743),
            .I(N__36738));
    InMux I__7684 (
            .O(N__36742),
            .I(N__36733));
    InMux I__7683 (
            .O(N__36741),
            .I(N__36733));
    LocalMux I__7682 (
            .O(N__36738),
            .I(measured_delay_hc_19));
    LocalMux I__7681 (
            .O(N__36733),
            .I(measured_delay_hc_19));
    CascadeMux I__7680 (
            .O(N__36728),
            .I(N__36725));
    InMux I__7679 (
            .O(N__36725),
            .I(N__36720));
    InMux I__7678 (
            .O(N__36724),
            .I(N__36717));
    InMux I__7677 (
            .O(N__36723),
            .I(N__36714));
    LocalMux I__7676 (
            .O(N__36720),
            .I(N__36709));
    LocalMux I__7675 (
            .O(N__36717),
            .I(N__36709));
    LocalMux I__7674 (
            .O(N__36714),
            .I(measured_delay_hc_22));
    Odrv4 I__7673 (
            .O(N__36709),
            .I(measured_delay_hc_22));
    InMux I__7672 (
            .O(N__36704),
            .I(N__36701));
    LocalMux I__7671 (
            .O(N__36701),
            .I(N__36693));
    InMux I__7670 (
            .O(N__36700),
            .I(N__36686));
    InMux I__7669 (
            .O(N__36699),
            .I(N__36686));
    InMux I__7668 (
            .O(N__36698),
            .I(N__36686));
    InMux I__7667 (
            .O(N__36697),
            .I(N__36681));
    InMux I__7666 (
            .O(N__36696),
            .I(N__36681));
    Span4Mux_v I__7665 (
            .O(N__36693),
            .I(N__36676));
    LocalMux I__7664 (
            .O(N__36686),
            .I(N__36676));
    LocalMux I__7663 (
            .O(N__36681),
            .I(N__36673));
    Span4Mux_h I__7662 (
            .O(N__36676),
            .I(N__36670));
    Span4Mux_v I__7661 (
            .O(N__36673),
            .I(N__36667));
    Span4Mux_v I__7660 (
            .O(N__36670),
            .I(N__36664));
    Span4Mux_h I__7659 (
            .O(N__36667),
            .I(N__36661));
    Span4Mux_h I__7658 (
            .O(N__36664),
            .I(N__36658));
    Span4Mux_h I__7657 (
            .O(N__36661),
            .I(N__36655));
    Odrv4 I__7656 (
            .O(N__36658),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    Odrv4 I__7655 (
            .O(N__36655),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    CascadeMux I__7654 (
            .O(N__36650),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_ ));
    InMux I__7653 (
            .O(N__36647),
            .I(N__36642));
    InMux I__7652 (
            .O(N__36646),
            .I(N__36637));
    InMux I__7651 (
            .O(N__36645),
            .I(N__36637));
    LocalMux I__7650 (
            .O(N__36642),
            .I(N__36634));
    LocalMux I__7649 (
            .O(N__36637),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__7648 (
            .O(N__36634),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__7647 (
            .O(N__36629),
            .I(N__36626));
    LocalMux I__7646 (
            .O(N__36626),
            .I(N__36623));
    Odrv4 I__7645 (
            .O(N__36623),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ));
    InMux I__7644 (
            .O(N__36620),
            .I(N__36617));
    LocalMux I__7643 (
            .O(N__36617),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12 ));
    InMux I__7642 (
            .O(N__36614),
            .I(N__36611));
    LocalMux I__7641 (
            .O(N__36611),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ));
    InMux I__7640 (
            .O(N__36608),
            .I(N__36605));
    LocalMux I__7639 (
            .O(N__36605),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0 ));
    CascadeMux I__7638 (
            .O(N__36602),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3_cascade_ ));
    InMux I__7637 (
            .O(N__36599),
            .I(N__36593));
    InMux I__7636 (
            .O(N__36598),
            .I(N__36590));
    InMux I__7635 (
            .O(N__36597),
            .I(N__36585));
    InMux I__7634 (
            .O(N__36596),
            .I(N__36585));
    LocalMux I__7633 (
            .O(N__36593),
            .I(N__36582));
    LocalMux I__7632 (
            .O(N__36590),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__7631 (
            .O(N__36585),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__7630 (
            .O(N__36582),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__7629 (
            .O(N__36575),
            .I(N__36570));
    InMux I__7628 (
            .O(N__36574),
            .I(N__36567));
    InMux I__7627 (
            .O(N__36573),
            .I(N__36564));
    LocalMux I__7626 (
            .O(N__36570),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__7625 (
            .O(N__36567),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__7624 (
            .O(N__36564),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    InMux I__7623 (
            .O(N__36557),
            .I(N__36554));
    LocalMux I__7622 (
            .O(N__36554),
            .I(N__36549));
    InMux I__7621 (
            .O(N__36553),
            .I(N__36546));
    InMux I__7620 (
            .O(N__36552),
            .I(N__36543));
    Odrv4 I__7619 (
            .O(N__36549),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__7618 (
            .O(N__36546),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__7617 (
            .O(N__36543),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__7616 (
            .O(N__36536),
            .I(N__36531));
    InMux I__7615 (
            .O(N__36535),
            .I(N__36526));
    InMux I__7614 (
            .O(N__36534),
            .I(N__36526));
    LocalMux I__7613 (
            .O(N__36531),
            .I(N__36520));
    LocalMux I__7612 (
            .O(N__36526),
            .I(N__36520));
    InMux I__7611 (
            .O(N__36525),
            .I(N__36517));
    Odrv4 I__7610 (
            .O(N__36520),
            .I(delay_tr_d2));
    LocalMux I__7609 (
            .O(N__36517),
            .I(delay_tr_d2));
    InMux I__7608 (
            .O(N__36512),
            .I(N__36509));
    LocalMux I__7607 (
            .O(N__36509),
            .I(N__36504));
    InMux I__7606 (
            .O(N__36508),
            .I(N__36501));
    InMux I__7605 (
            .O(N__36507),
            .I(N__36498));
    Odrv4 I__7604 (
            .O(N__36504),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__7603 (
            .O(N__36501),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__7602 (
            .O(N__36498),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__7601 (
            .O(N__36491),
            .I(N__36486));
    InMux I__7600 (
            .O(N__36490),
            .I(N__36483));
    InMux I__7599 (
            .O(N__36489),
            .I(N__36480));
    LocalMux I__7598 (
            .O(N__36486),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__7597 (
            .O(N__36483),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__7596 (
            .O(N__36480),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__7595 (
            .O(N__36473),
            .I(N__36470));
    LocalMux I__7594 (
            .O(N__36470),
            .I(N__36467));
    Span4Mux_h I__7593 (
            .O(N__36467),
            .I(N__36464));
    Sp12to4 I__7592 (
            .O(N__36464),
            .I(N__36461));
    Odrv12 I__7591 (
            .O(N__36461),
            .I(delay_hc_input_c));
    InMux I__7590 (
            .O(N__36458),
            .I(N__36455));
    LocalMux I__7589 (
            .O(N__36455),
            .I(delay_hc_d1));
    InMux I__7588 (
            .O(N__36452),
            .I(N__36448));
    InMux I__7587 (
            .O(N__36451),
            .I(N__36445));
    LocalMux I__7586 (
            .O(N__36448),
            .I(N__36442));
    LocalMux I__7585 (
            .O(N__36445),
            .I(N__36437));
    Span4Mux_h I__7584 (
            .O(N__36442),
            .I(N__36434));
    InMux I__7583 (
            .O(N__36441),
            .I(N__36431));
    InMux I__7582 (
            .O(N__36440),
            .I(N__36428));
    Odrv4 I__7581 (
            .O(N__36437),
            .I(delay_hc_d2));
    Odrv4 I__7580 (
            .O(N__36434),
            .I(delay_hc_d2));
    LocalMux I__7579 (
            .O(N__36431),
            .I(delay_hc_d2));
    LocalMux I__7578 (
            .O(N__36428),
            .I(delay_hc_d2));
    CascadeMux I__7577 (
            .O(N__36419),
            .I(N__36414));
    InMux I__7576 (
            .O(N__36418),
            .I(N__36410));
    InMux I__7575 (
            .O(N__36417),
            .I(N__36407));
    InMux I__7574 (
            .O(N__36414),
            .I(N__36404));
    CascadeMux I__7573 (
            .O(N__36413),
            .I(N__36400));
    LocalMux I__7572 (
            .O(N__36410),
            .I(N__36397));
    LocalMux I__7571 (
            .O(N__36407),
            .I(N__36394));
    LocalMux I__7570 (
            .O(N__36404),
            .I(N__36391));
    InMux I__7569 (
            .O(N__36403),
            .I(N__36388));
    InMux I__7568 (
            .O(N__36400),
            .I(N__36385));
    Span12Mux_s11_h I__7567 (
            .O(N__36397),
            .I(N__36382));
    Sp12to4 I__7566 (
            .O(N__36394),
            .I(N__36379));
    Span4Mux_v I__7565 (
            .O(N__36391),
            .I(N__36374));
    LocalMux I__7564 (
            .O(N__36388),
            .I(N__36374));
    LocalMux I__7563 (
            .O(N__36385),
            .I(measured_delay_hc_9));
    Odrv12 I__7562 (
            .O(N__36382),
            .I(measured_delay_hc_9));
    Odrv12 I__7561 (
            .O(N__36379),
            .I(measured_delay_hc_9));
    Odrv4 I__7560 (
            .O(N__36374),
            .I(measured_delay_hc_9));
    InMux I__7559 (
            .O(N__36365),
            .I(N__36361));
    InMux I__7558 (
            .O(N__36364),
            .I(N__36358));
    LocalMux I__7557 (
            .O(N__36361),
            .I(N__36353));
    LocalMux I__7556 (
            .O(N__36358),
            .I(N__36353));
    Odrv4 I__7555 (
            .O(N__36353),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__7554 (
            .O(N__36350),
            .I(N__36347));
    LocalMux I__7553 (
            .O(N__36347),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__7552 (
            .O(N__36344),
            .I(N__36341));
    LocalMux I__7551 (
            .O(N__36341),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__7550 (
            .O(N__36338),
            .I(N__36335));
    LocalMux I__7549 (
            .O(N__36335),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__7548 (
            .O(N__36332),
            .I(N__36329));
    LocalMux I__7547 (
            .O(N__36329),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__7546 (
            .O(N__36326),
            .I(N__36312));
    InMux I__7545 (
            .O(N__36325),
            .I(N__36295));
    InMux I__7544 (
            .O(N__36324),
            .I(N__36295));
    InMux I__7543 (
            .O(N__36323),
            .I(N__36295));
    InMux I__7542 (
            .O(N__36322),
            .I(N__36295));
    InMux I__7541 (
            .O(N__36321),
            .I(N__36295));
    InMux I__7540 (
            .O(N__36320),
            .I(N__36295));
    InMux I__7539 (
            .O(N__36319),
            .I(N__36295));
    InMux I__7538 (
            .O(N__36318),
            .I(N__36295));
    InMux I__7537 (
            .O(N__36317),
            .I(N__36280));
    InMux I__7536 (
            .O(N__36316),
            .I(N__36280));
    InMux I__7535 (
            .O(N__36315),
            .I(N__36280));
    LocalMux I__7534 (
            .O(N__36312),
            .I(N__36273));
    LocalMux I__7533 (
            .O(N__36295),
            .I(N__36273));
    InMux I__7532 (
            .O(N__36294),
            .I(N__36256));
    InMux I__7531 (
            .O(N__36293),
            .I(N__36256));
    InMux I__7530 (
            .O(N__36292),
            .I(N__36256));
    InMux I__7529 (
            .O(N__36291),
            .I(N__36256));
    InMux I__7528 (
            .O(N__36290),
            .I(N__36256));
    InMux I__7527 (
            .O(N__36289),
            .I(N__36256));
    InMux I__7526 (
            .O(N__36288),
            .I(N__36256));
    InMux I__7525 (
            .O(N__36287),
            .I(N__36256));
    LocalMux I__7524 (
            .O(N__36280),
            .I(N__36252));
    InMux I__7523 (
            .O(N__36279),
            .I(N__36249));
    InMux I__7522 (
            .O(N__36278),
            .I(N__36246));
    Span4Mux_v I__7521 (
            .O(N__36273),
            .I(N__36240));
    LocalMux I__7520 (
            .O(N__36256),
            .I(N__36240));
    InMux I__7519 (
            .O(N__36255),
            .I(N__36237));
    Span4Mux_h I__7518 (
            .O(N__36252),
            .I(N__36232));
    LocalMux I__7517 (
            .O(N__36249),
            .I(N__36232));
    LocalMux I__7516 (
            .O(N__36246),
            .I(N__36229));
    InMux I__7515 (
            .O(N__36245),
            .I(N__36226));
    Span4Mux_v I__7514 (
            .O(N__36240),
            .I(N__36223));
    LocalMux I__7513 (
            .O(N__36237),
            .I(N__36216));
    Sp12to4 I__7512 (
            .O(N__36232),
            .I(N__36216));
    Sp12to4 I__7511 (
            .O(N__36229),
            .I(N__36216));
    LocalMux I__7510 (
            .O(N__36226),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__7509 (
            .O(N__36223),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv12 I__7508 (
            .O(N__36216),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__7507 (
            .O(N__36209),
            .I(N__36201));
    CascadeMux I__7506 (
            .O(N__36208),
            .I(N__36198));
    CascadeMux I__7505 (
            .O(N__36207),
            .I(N__36194));
    CascadeMux I__7504 (
            .O(N__36206),
            .I(N__36188));
    CascadeMux I__7503 (
            .O(N__36205),
            .I(N__36185));
    CascadeMux I__7502 (
            .O(N__36204),
            .I(N__36177));
    InMux I__7501 (
            .O(N__36201),
            .I(N__36173));
    InMux I__7500 (
            .O(N__36198),
            .I(N__36156));
    InMux I__7499 (
            .O(N__36197),
            .I(N__36156));
    InMux I__7498 (
            .O(N__36194),
            .I(N__36156));
    InMux I__7497 (
            .O(N__36193),
            .I(N__36156));
    InMux I__7496 (
            .O(N__36192),
            .I(N__36156));
    InMux I__7495 (
            .O(N__36191),
            .I(N__36156));
    InMux I__7494 (
            .O(N__36188),
            .I(N__36156));
    InMux I__7493 (
            .O(N__36185),
            .I(N__36156));
    CascadeMux I__7492 (
            .O(N__36184),
            .I(N__36152));
    CascadeMux I__7491 (
            .O(N__36183),
            .I(N__36149));
    CascadeMux I__7490 (
            .O(N__36182),
            .I(N__36145));
    CascadeMux I__7489 (
            .O(N__36181),
            .I(N__36140));
    CascadeMux I__7488 (
            .O(N__36180),
            .I(N__36137));
    InMux I__7487 (
            .O(N__36177),
            .I(N__36134));
    CascadeMux I__7486 (
            .O(N__36176),
            .I(N__36131));
    LocalMux I__7485 (
            .O(N__36173),
            .I(N__36126));
    LocalMux I__7484 (
            .O(N__36156),
            .I(N__36126));
    InMux I__7483 (
            .O(N__36155),
            .I(N__36109));
    InMux I__7482 (
            .O(N__36152),
            .I(N__36109));
    InMux I__7481 (
            .O(N__36149),
            .I(N__36109));
    InMux I__7480 (
            .O(N__36148),
            .I(N__36109));
    InMux I__7479 (
            .O(N__36145),
            .I(N__36109));
    InMux I__7478 (
            .O(N__36144),
            .I(N__36109));
    InMux I__7477 (
            .O(N__36143),
            .I(N__36109));
    InMux I__7476 (
            .O(N__36140),
            .I(N__36109));
    InMux I__7475 (
            .O(N__36137),
            .I(N__36106));
    LocalMux I__7474 (
            .O(N__36134),
            .I(N__36099));
    InMux I__7473 (
            .O(N__36131),
            .I(N__36096));
    Span4Mux_v I__7472 (
            .O(N__36126),
            .I(N__36091));
    LocalMux I__7471 (
            .O(N__36109),
            .I(N__36091));
    LocalMux I__7470 (
            .O(N__36106),
            .I(N__36088));
    InMux I__7469 (
            .O(N__36105),
            .I(N__36081));
    InMux I__7468 (
            .O(N__36104),
            .I(N__36081));
    InMux I__7467 (
            .O(N__36103),
            .I(N__36081));
    InMux I__7466 (
            .O(N__36102),
            .I(N__36078));
    Odrv12 I__7465 (
            .O(N__36099),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__7464 (
            .O(N__36096),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__7463 (
            .O(N__36091),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__7462 (
            .O(N__36088),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__7461 (
            .O(N__36081),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__7460 (
            .O(N__36078),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__7459 (
            .O(N__36065),
            .I(N__36057));
    CascadeMux I__7458 (
            .O(N__36064),
            .I(N__36047));
    CascadeMux I__7457 (
            .O(N__36063),
            .I(N__36044));
    CascadeMux I__7456 (
            .O(N__36062),
            .I(N__36041));
    CascadeMux I__7455 (
            .O(N__36061),
            .I(N__36038));
    InMux I__7454 (
            .O(N__36060),
            .I(N__36031));
    LocalMux I__7453 (
            .O(N__36057),
            .I(N__36028));
    CascadeMux I__7452 (
            .O(N__36056),
            .I(N__36025));
    CascadeMux I__7451 (
            .O(N__36055),
            .I(N__36022));
    InMux I__7450 (
            .O(N__36054),
            .I(N__36018));
    CascadeMux I__7449 (
            .O(N__36053),
            .I(N__36013));
    CascadeMux I__7448 (
            .O(N__36052),
            .I(N__36010));
    CascadeMux I__7447 (
            .O(N__36051),
            .I(N__36007));
    CascadeMux I__7446 (
            .O(N__36050),
            .I(N__36004));
    InMux I__7445 (
            .O(N__36047),
            .I(N__35991));
    InMux I__7444 (
            .O(N__36044),
            .I(N__35991));
    InMux I__7443 (
            .O(N__36041),
            .I(N__35991));
    InMux I__7442 (
            .O(N__36038),
            .I(N__35991));
    InMux I__7441 (
            .O(N__36037),
            .I(N__35982));
    InMux I__7440 (
            .O(N__36036),
            .I(N__35982));
    InMux I__7439 (
            .O(N__36035),
            .I(N__35982));
    InMux I__7438 (
            .O(N__36034),
            .I(N__35982));
    LocalMux I__7437 (
            .O(N__36031),
            .I(N__35979));
    Span4Mux_v I__7436 (
            .O(N__36028),
            .I(N__35976));
    InMux I__7435 (
            .O(N__36025),
            .I(N__35969));
    InMux I__7434 (
            .O(N__36022),
            .I(N__35969));
    InMux I__7433 (
            .O(N__36021),
            .I(N__35969));
    LocalMux I__7432 (
            .O(N__36018),
            .I(N__35966));
    InMux I__7431 (
            .O(N__36017),
            .I(N__35963));
    InMux I__7430 (
            .O(N__36016),
            .I(N__35960));
    InMux I__7429 (
            .O(N__36013),
            .I(N__35951));
    InMux I__7428 (
            .O(N__36010),
            .I(N__35951));
    InMux I__7427 (
            .O(N__36007),
            .I(N__35951));
    InMux I__7426 (
            .O(N__36004),
            .I(N__35951));
    InMux I__7425 (
            .O(N__36003),
            .I(N__35942));
    InMux I__7424 (
            .O(N__36002),
            .I(N__35942));
    InMux I__7423 (
            .O(N__36001),
            .I(N__35942));
    InMux I__7422 (
            .O(N__36000),
            .I(N__35942));
    LocalMux I__7421 (
            .O(N__35991),
            .I(N__35933));
    LocalMux I__7420 (
            .O(N__35982),
            .I(N__35933));
    Span4Mux_h I__7419 (
            .O(N__35979),
            .I(N__35933));
    Span4Mux_v I__7418 (
            .O(N__35976),
            .I(N__35933));
    LocalMux I__7417 (
            .O(N__35969),
            .I(N__35930));
    Span4Mux_v I__7416 (
            .O(N__35966),
            .I(N__35925));
    LocalMux I__7415 (
            .O(N__35963),
            .I(N__35925));
    LocalMux I__7414 (
            .O(N__35960),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__7413 (
            .O(N__35951),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__7412 (
            .O(N__35942),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__7411 (
            .O(N__35933),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__7410 (
            .O(N__35930),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__7409 (
            .O(N__35925),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__7408 (
            .O(N__35912),
            .I(N__35909));
    LocalMux I__7407 (
            .O(N__35909),
            .I(N__35906));
    Odrv12 I__7406 (
            .O(N__35906),
            .I(delay_tr_input_c));
    InMux I__7405 (
            .O(N__35903),
            .I(N__35900));
    LocalMux I__7404 (
            .O(N__35900),
            .I(delay_tr_d1));
    CEMux I__7403 (
            .O(N__35897),
            .I(N__35894));
    LocalMux I__7402 (
            .O(N__35894),
            .I(N__35891));
    Span4Mux_h I__7401 (
            .O(N__35891),
            .I(N__35888));
    Span4Mux_v I__7400 (
            .O(N__35888),
            .I(N__35884));
    CEMux I__7399 (
            .O(N__35887),
            .I(N__35881));
    Span4Mux_v I__7398 (
            .O(N__35884),
            .I(N__35874));
    LocalMux I__7397 (
            .O(N__35881),
            .I(N__35874));
    IoInMux I__7396 (
            .O(N__35880),
            .I(N__35871));
    CEMux I__7395 (
            .O(N__35879),
            .I(N__35868));
    Span4Mux_v I__7394 (
            .O(N__35874),
            .I(N__35865));
    LocalMux I__7393 (
            .O(N__35871),
            .I(N__35862));
    LocalMux I__7392 (
            .O(N__35868),
            .I(N__35858));
    Span4Mux_v I__7391 (
            .O(N__35865),
            .I(N__35855));
    IoSpan4Mux I__7390 (
            .O(N__35862),
            .I(N__35852));
    CEMux I__7389 (
            .O(N__35861),
            .I(N__35849));
    Span12Mux_h I__7388 (
            .O(N__35858),
            .I(N__35846));
    Span4Mux_v I__7387 (
            .O(N__35855),
            .I(N__35841));
    Span4Mux_s0_v I__7386 (
            .O(N__35852),
            .I(N__35841));
    LocalMux I__7385 (
            .O(N__35849),
            .I(N__35838));
    Span12Mux_v I__7384 (
            .O(N__35846),
            .I(N__35833));
    Span4Mux_v I__7383 (
            .O(N__35841),
            .I(N__35828));
    Span4Mux_h I__7382 (
            .O(N__35838),
            .I(N__35828));
    CEMux I__7381 (
            .O(N__35837),
            .I(N__35825));
    CEMux I__7380 (
            .O(N__35836),
            .I(N__35822));
    Odrv12 I__7379 (
            .O(N__35833),
            .I(red_c_i));
    Odrv4 I__7378 (
            .O(N__35828),
            .I(red_c_i));
    LocalMux I__7377 (
            .O(N__35825),
            .I(red_c_i));
    LocalMux I__7376 (
            .O(N__35822),
            .I(red_c_i));
    InMux I__7375 (
            .O(N__35813),
            .I(N__35810));
    LocalMux I__7374 (
            .O(N__35810),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__7373 (
            .O(N__35807),
            .I(N__35804));
    LocalMux I__7372 (
            .O(N__35804),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__7371 (
            .O(N__35801),
            .I(N__35798));
    LocalMux I__7370 (
            .O(N__35798),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__7369 (
            .O(N__35795),
            .I(N__35792));
    LocalMux I__7368 (
            .O(N__35792),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__7367 (
            .O(N__35789),
            .I(N__35786));
    LocalMux I__7366 (
            .O(N__35786),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__7365 (
            .O(N__35783),
            .I(N__35780));
    LocalMux I__7364 (
            .O(N__35780),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__7363 (
            .O(N__35777),
            .I(N__35774));
    LocalMux I__7362 (
            .O(N__35774),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__7361 (
            .O(N__35771),
            .I(N__35768));
    LocalMux I__7360 (
            .O(N__35768),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__7359 (
            .O(N__35765),
            .I(N__35762));
    LocalMux I__7358 (
            .O(N__35762),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__7357 (
            .O(N__35759),
            .I(N__35756));
    LocalMux I__7356 (
            .O(N__35756),
            .I(N__35753));
    Odrv4 I__7355 (
            .O(N__35753),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__7354 (
            .O(N__35750),
            .I(N__35747));
    LocalMux I__7353 (
            .O(N__35747),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__7352 (
            .O(N__35744),
            .I(N__35741));
    LocalMux I__7351 (
            .O(N__35741),
            .I(N__35738));
    Odrv4 I__7350 (
            .O(N__35738),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__7349 (
            .O(N__35735),
            .I(N__35732));
    LocalMux I__7348 (
            .O(N__35732),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__7347 (
            .O(N__35729),
            .I(N__35726));
    LocalMux I__7346 (
            .O(N__35726),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__7345 (
            .O(N__35723),
            .I(N__35720));
    LocalMux I__7344 (
            .O(N__35720),
            .I(N__35717));
    Span12Mux_s9_v I__7343 (
            .O(N__35717),
            .I(N__35714));
    Odrv12 I__7342 (
            .O(N__35714),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ));
    InMux I__7341 (
            .O(N__35711),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__7340 (
            .O(N__35708),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__7339 (
            .O(N__35705),
            .I(N__35702));
    LocalMux I__7338 (
            .O(N__35702),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__7337 (
            .O(N__35699),
            .I(N__35696));
    LocalMux I__7336 (
            .O(N__35696),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__7335 (
            .O(N__35693),
            .I(N__35690));
    LocalMux I__7334 (
            .O(N__35690),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__7333 (
            .O(N__35687),
            .I(N__35684));
    LocalMux I__7332 (
            .O(N__35684),
            .I(N__35681));
    Odrv12 I__7331 (
            .O(N__35681),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__7330 (
            .O(N__35678),
            .I(N__35675));
    LocalMux I__7329 (
            .O(N__35675),
            .I(N__35672));
    Odrv4 I__7328 (
            .O(N__35672),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__7327 (
            .O(N__35669),
            .I(N__35666));
    LocalMux I__7326 (
            .O(N__35666),
            .I(N__35663));
    Odrv4 I__7325 (
            .O(N__35663),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__7324 (
            .O(N__35660),
            .I(N__35657));
    LocalMux I__7323 (
            .O(N__35657),
            .I(N__35654));
    Odrv4 I__7322 (
            .O(N__35654),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__7321 (
            .O(N__35651),
            .I(bfn_14_19_0_));
    InMux I__7320 (
            .O(N__35648),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__7319 (
            .O(N__35645),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__7318 (
            .O(N__35642),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__7317 (
            .O(N__35639),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__7316 (
            .O(N__35636),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__7315 (
            .O(N__35633),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__7314 (
            .O(N__35630),
            .I(N__35627));
    LocalMux I__7313 (
            .O(N__35627),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__7312 (
            .O(N__35624),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__7311 (
            .O(N__35621),
            .I(bfn_14_20_0_));
    CascadeMux I__7310 (
            .O(N__35618),
            .I(N__35612));
    InMux I__7309 (
            .O(N__35617),
            .I(N__35605));
    InMux I__7308 (
            .O(N__35616),
            .I(N__35605));
    CascadeMux I__7307 (
            .O(N__35615),
            .I(N__35601));
    InMux I__7306 (
            .O(N__35612),
            .I(N__35587));
    InMux I__7305 (
            .O(N__35611),
            .I(N__35587));
    InMux I__7304 (
            .O(N__35610),
            .I(N__35587));
    LocalMux I__7303 (
            .O(N__35605),
            .I(N__35580));
    InMux I__7302 (
            .O(N__35604),
            .I(N__35577));
    InMux I__7301 (
            .O(N__35601),
            .I(N__35568));
    InMux I__7300 (
            .O(N__35600),
            .I(N__35568));
    InMux I__7299 (
            .O(N__35599),
            .I(N__35568));
    InMux I__7298 (
            .O(N__35598),
            .I(N__35568));
    InMux I__7297 (
            .O(N__35597),
            .I(N__35559));
    InMux I__7296 (
            .O(N__35596),
            .I(N__35559));
    InMux I__7295 (
            .O(N__35595),
            .I(N__35559));
    InMux I__7294 (
            .O(N__35594),
            .I(N__35559));
    LocalMux I__7293 (
            .O(N__35587),
            .I(N__35556));
    InMux I__7292 (
            .O(N__35586),
            .I(N__35547));
    InMux I__7291 (
            .O(N__35585),
            .I(N__35547));
    InMux I__7290 (
            .O(N__35584),
            .I(N__35547));
    InMux I__7289 (
            .O(N__35583),
            .I(N__35547));
    Span4Mux_h I__7288 (
            .O(N__35580),
            .I(N__35544));
    LocalMux I__7287 (
            .O(N__35577),
            .I(N__35537));
    LocalMux I__7286 (
            .O(N__35568),
            .I(N__35528));
    LocalMux I__7285 (
            .O(N__35559),
            .I(N__35528));
    Span4Mux_v I__7284 (
            .O(N__35556),
            .I(N__35528));
    LocalMux I__7283 (
            .O(N__35547),
            .I(N__35528));
    Span4Mux_h I__7282 (
            .O(N__35544),
            .I(N__35525));
    InMux I__7281 (
            .O(N__35543),
            .I(N__35516));
    InMux I__7280 (
            .O(N__35542),
            .I(N__35516));
    InMux I__7279 (
            .O(N__35541),
            .I(N__35516));
    InMux I__7278 (
            .O(N__35540),
            .I(N__35516));
    Span4Mux_h I__7277 (
            .O(N__35537),
            .I(N__35513));
    Span4Mux_v I__7276 (
            .O(N__35528),
            .I(N__35508));
    Span4Mux_h I__7275 (
            .O(N__35525),
            .I(N__35508));
    LocalMux I__7274 (
            .O(N__35516),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__7273 (
            .O(N__35513),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__7272 (
            .O(N__35508),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    InMux I__7271 (
            .O(N__35501),
            .I(N__35496));
    CascadeMux I__7270 (
            .O(N__35500),
            .I(N__35493));
    InMux I__7269 (
            .O(N__35499),
            .I(N__35490));
    LocalMux I__7268 (
            .O(N__35496),
            .I(N__35485));
    InMux I__7267 (
            .O(N__35493),
            .I(N__35482));
    LocalMux I__7266 (
            .O(N__35490),
            .I(N__35479));
    InMux I__7265 (
            .O(N__35489),
            .I(N__35476));
    InMux I__7264 (
            .O(N__35488),
            .I(N__35473));
    Span4Mux_v I__7263 (
            .O(N__35485),
            .I(N__35470));
    LocalMux I__7262 (
            .O(N__35482),
            .I(N__35467));
    Span4Mux_v I__7261 (
            .O(N__35479),
            .I(N__35462));
    LocalMux I__7260 (
            .O(N__35476),
            .I(N__35462));
    LocalMux I__7259 (
            .O(N__35473),
            .I(measured_delay_hc_8));
    Odrv4 I__7258 (
            .O(N__35470),
            .I(measured_delay_hc_8));
    Odrv12 I__7257 (
            .O(N__35467),
            .I(measured_delay_hc_8));
    Odrv4 I__7256 (
            .O(N__35462),
            .I(measured_delay_hc_8));
    InMux I__7255 (
            .O(N__35453),
            .I(N__35440));
    InMux I__7254 (
            .O(N__35452),
            .I(N__35440));
    InMux I__7253 (
            .O(N__35451),
            .I(N__35440));
    InMux I__7252 (
            .O(N__35450),
            .I(N__35427));
    InMux I__7251 (
            .O(N__35449),
            .I(N__35427));
    InMux I__7250 (
            .O(N__35448),
            .I(N__35427));
    InMux I__7249 (
            .O(N__35447),
            .I(N__35427));
    LocalMux I__7248 (
            .O(N__35440),
            .I(N__35424));
    InMux I__7247 (
            .O(N__35439),
            .I(N__35415));
    InMux I__7246 (
            .O(N__35438),
            .I(N__35415));
    InMux I__7245 (
            .O(N__35437),
            .I(N__35415));
    InMux I__7244 (
            .O(N__35436),
            .I(N__35415));
    LocalMux I__7243 (
            .O(N__35427),
            .I(N__35409));
    Span4Mux_v I__7242 (
            .O(N__35424),
            .I(N__35404));
    LocalMux I__7241 (
            .O(N__35415),
            .I(N__35404));
    InMux I__7240 (
            .O(N__35414),
            .I(N__35397));
    InMux I__7239 (
            .O(N__35413),
            .I(N__35397));
    InMux I__7238 (
            .O(N__35412),
            .I(N__35397));
    Odrv12 I__7237 (
            .O(N__35409),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    Odrv4 I__7236 (
            .O(N__35404),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    LocalMux I__7235 (
            .O(N__35397),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    InMux I__7234 (
            .O(N__35390),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__7233 (
            .O(N__35387),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__7232 (
            .O(N__35384),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__7231 (
            .O(N__35381),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__7230 (
            .O(N__35378),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__7229 (
            .O(N__35375),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__7228 (
            .O(N__35372),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__7227 (
            .O(N__35369),
            .I(N__35365));
    CascadeMux I__7226 (
            .O(N__35368),
            .I(N__35361));
    LocalMux I__7225 (
            .O(N__35365),
            .I(N__35357));
    InMux I__7224 (
            .O(N__35364),
            .I(N__35354));
    InMux I__7223 (
            .O(N__35361),
            .I(N__35351));
    CascadeMux I__7222 (
            .O(N__35360),
            .I(N__35347));
    Sp12to4 I__7221 (
            .O(N__35357),
            .I(N__35342));
    LocalMux I__7220 (
            .O(N__35354),
            .I(N__35342));
    LocalMux I__7219 (
            .O(N__35351),
            .I(N__35339));
    CascadeMux I__7218 (
            .O(N__35350),
            .I(N__35336));
    InMux I__7217 (
            .O(N__35347),
            .I(N__35333));
    Span12Mux_v I__7216 (
            .O(N__35342),
            .I(N__35330));
    Span4Mux_h I__7215 (
            .O(N__35339),
            .I(N__35327));
    InMux I__7214 (
            .O(N__35336),
            .I(N__35324));
    LocalMux I__7213 (
            .O(N__35333),
            .I(measured_delay_hc_12));
    Odrv12 I__7212 (
            .O(N__35330),
            .I(measured_delay_hc_12));
    Odrv4 I__7211 (
            .O(N__35327),
            .I(measured_delay_hc_12));
    LocalMux I__7210 (
            .O(N__35324),
            .I(measured_delay_hc_12));
    InMux I__7209 (
            .O(N__35315),
            .I(N__35312));
    LocalMux I__7208 (
            .O(N__35312),
            .I(N__35308));
    InMux I__7207 (
            .O(N__35311),
            .I(N__35305));
    Span4Mux_v I__7206 (
            .O(N__35308),
            .I(N__35298));
    LocalMux I__7205 (
            .O(N__35305),
            .I(N__35298));
    InMux I__7204 (
            .O(N__35304),
            .I(N__35295));
    InMux I__7203 (
            .O(N__35303),
            .I(N__35292));
    Span4Mux_h I__7202 (
            .O(N__35298),
            .I(N__35289));
    LocalMux I__7201 (
            .O(N__35295),
            .I(N__35286));
    LocalMux I__7200 (
            .O(N__35292),
            .I(measured_delay_hc_1));
    Odrv4 I__7199 (
            .O(N__35289),
            .I(measured_delay_hc_1));
    Odrv12 I__7198 (
            .O(N__35286),
            .I(measured_delay_hc_1));
    CascadeMux I__7197 (
            .O(N__35279),
            .I(N__35275));
    CascadeMux I__7196 (
            .O(N__35278),
            .I(N__35271));
    InMux I__7195 (
            .O(N__35275),
            .I(N__35268));
    CascadeMux I__7194 (
            .O(N__35274),
            .I(N__35264));
    InMux I__7193 (
            .O(N__35271),
            .I(N__35261));
    LocalMux I__7192 (
            .O(N__35268),
            .I(N__35258));
    InMux I__7191 (
            .O(N__35267),
            .I(N__35253));
    InMux I__7190 (
            .O(N__35264),
            .I(N__35253));
    LocalMux I__7189 (
            .O(N__35261),
            .I(N__35249));
    Span4Mux_v I__7188 (
            .O(N__35258),
            .I(N__35244));
    LocalMux I__7187 (
            .O(N__35253),
            .I(N__35244));
    InMux I__7186 (
            .O(N__35252),
            .I(N__35241));
    Span12Mux_h I__7185 (
            .O(N__35249),
            .I(N__35238));
    Span4Mux_v I__7184 (
            .O(N__35244),
            .I(N__35235));
    LocalMux I__7183 (
            .O(N__35241),
            .I(measured_delay_hc_3));
    Odrv12 I__7182 (
            .O(N__35238),
            .I(measured_delay_hc_3));
    Odrv4 I__7181 (
            .O(N__35235),
            .I(measured_delay_hc_3));
    InMux I__7180 (
            .O(N__35228),
            .I(N__35225));
    LocalMux I__7179 (
            .O(N__35225),
            .I(N__35222));
    Span4Mux_h I__7178 (
            .O(N__35222),
            .I(N__35218));
    InMux I__7177 (
            .O(N__35221),
            .I(N__35215));
    Span4Mux_v I__7176 (
            .O(N__35218),
            .I(N__35210));
    LocalMux I__7175 (
            .O(N__35215),
            .I(N__35207));
    InMux I__7174 (
            .O(N__35214),
            .I(N__35202));
    InMux I__7173 (
            .O(N__35213),
            .I(N__35202));
    Odrv4 I__7172 (
            .O(N__35210),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    Odrv12 I__7171 (
            .O(N__35207),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    LocalMux I__7170 (
            .O(N__35202),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    InMux I__7169 (
            .O(N__35195),
            .I(N__35191));
    CascadeMux I__7168 (
            .O(N__35194),
            .I(N__35188));
    LocalMux I__7167 (
            .O(N__35191),
            .I(N__35184));
    InMux I__7166 (
            .O(N__35188),
            .I(N__35181));
    InMux I__7165 (
            .O(N__35187),
            .I(N__35177));
    Span4Mux_v I__7164 (
            .O(N__35184),
            .I(N__35173));
    LocalMux I__7163 (
            .O(N__35181),
            .I(N__35170));
    InMux I__7162 (
            .O(N__35180),
            .I(N__35167));
    LocalMux I__7161 (
            .O(N__35177),
            .I(N__35164));
    InMux I__7160 (
            .O(N__35176),
            .I(N__35161));
    Span4Mux_v I__7159 (
            .O(N__35173),
            .I(N__35158));
    Span4Mux_v I__7158 (
            .O(N__35170),
            .I(N__35151));
    LocalMux I__7157 (
            .O(N__35167),
            .I(N__35151));
    Span4Mux_h I__7156 (
            .O(N__35164),
            .I(N__35151));
    LocalMux I__7155 (
            .O(N__35161),
            .I(measured_delay_hc_15));
    Odrv4 I__7154 (
            .O(N__35158),
            .I(measured_delay_hc_15));
    Odrv4 I__7153 (
            .O(N__35151),
            .I(measured_delay_hc_15));
    InMux I__7152 (
            .O(N__35144),
            .I(N__35140));
    InMux I__7151 (
            .O(N__35143),
            .I(N__35137));
    LocalMux I__7150 (
            .O(N__35140),
            .I(N__35133));
    LocalMux I__7149 (
            .O(N__35137),
            .I(N__35128));
    InMux I__7148 (
            .O(N__35136),
            .I(N__35125));
    Span4Mux_v I__7147 (
            .O(N__35133),
            .I(N__35122));
    InMux I__7146 (
            .O(N__35132),
            .I(N__35119));
    InMux I__7145 (
            .O(N__35131),
            .I(N__35116));
    Span12Mux_v I__7144 (
            .O(N__35128),
            .I(N__35113));
    LocalMux I__7143 (
            .O(N__35125),
            .I(N__35110));
    Span4Mux_v I__7142 (
            .O(N__35122),
            .I(N__35105));
    LocalMux I__7141 (
            .O(N__35119),
            .I(N__35105));
    LocalMux I__7140 (
            .O(N__35116),
            .I(measured_delay_hc_13));
    Odrv12 I__7139 (
            .O(N__35113),
            .I(measured_delay_hc_13));
    Odrv12 I__7138 (
            .O(N__35110),
            .I(measured_delay_hc_13));
    Odrv4 I__7137 (
            .O(N__35105),
            .I(measured_delay_hc_13));
    InMux I__7136 (
            .O(N__35096),
            .I(N__35092));
    CascadeMux I__7135 (
            .O(N__35095),
            .I(N__35086));
    LocalMux I__7134 (
            .O(N__35092),
            .I(N__35083));
    InMux I__7133 (
            .O(N__35091),
            .I(N__35080));
    InMux I__7132 (
            .O(N__35090),
            .I(N__35075));
    InMux I__7131 (
            .O(N__35089),
            .I(N__35075));
    InMux I__7130 (
            .O(N__35086),
            .I(N__35072));
    Sp12to4 I__7129 (
            .O(N__35083),
            .I(N__35067));
    LocalMux I__7128 (
            .O(N__35080),
            .I(N__35067));
    LocalMux I__7127 (
            .O(N__35075),
            .I(N__35064));
    LocalMux I__7126 (
            .O(N__35072),
            .I(measured_delay_hc_18));
    Odrv12 I__7125 (
            .O(N__35067),
            .I(measured_delay_hc_18));
    Odrv4 I__7124 (
            .O(N__35064),
            .I(measured_delay_hc_18));
    InMux I__7123 (
            .O(N__35057),
            .I(N__35053));
    InMux I__7122 (
            .O(N__35056),
            .I(N__35050));
    LocalMux I__7121 (
            .O(N__35053),
            .I(N__35047));
    LocalMux I__7120 (
            .O(N__35050),
            .I(N__35040));
    Span4Mux_h I__7119 (
            .O(N__35047),
            .I(N__35040));
    InMux I__7118 (
            .O(N__35046),
            .I(N__35036));
    InMux I__7117 (
            .O(N__35045),
            .I(N__35033));
    Span4Mux_v I__7116 (
            .O(N__35040),
            .I(N__35030));
    InMux I__7115 (
            .O(N__35039),
            .I(N__35027));
    LocalMux I__7114 (
            .O(N__35036),
            .I(N__35024));
    LocalMux I__7113 (
            .O(N__35033),
            .I(measured_delay_hc_6));
    Odrv4 I__7112 (
            .O(N__35030),
            .I(measured_delay_hc_6));
    LocalMux I__7111 (
            .O(N__35027),
            .I(measured_delay_hc_6));
    Odrv4 I__7110 (
            .O(N__35024),
            .I(measured_delay_hc_6));
    InMux I__7109 (
            .O(N__35015),
            .I(N__35002));
    InMux I__7108 (
            .O(N__35014),
            .I(N__35002));
    InMux I__7107 (
            .O(N__35013),
            .I(N__35002));
    InMux I__7106 (
            .O(N__35012),
            .I(N__34993));
    InMux I__7105 (
            .O(N__35011),
            .I(N__34993));
    InMux I__7104 (
            .O(N__35010),
            .I(N__34993));
    InMux I__7103 (
            .O(N__35009),
            .I(N__34993));
    LocalMux I__7102 (
            .O(N__35002),
            .I(N__34982));
    LocalMux I__7101 (
            .O(N__34993),
            .I(N__34979));
    InMux I__7100 (
            .O(N__34992),
            .I(N__34976));
    InMux I__7099 (
            .O(N__34991),
            .I(N__34969));
    InMux I__7098 (
            .O(N__34990),
            .I(N__34969));
    InMux I__7097 (
            .O(N__34989),
            .I(N__34969));
    InMux I__7096 (
            .O(N__34988),
            .I(N__34964));
    InMux I__7095 (
            .O(N__34987),
            .I(N__34964));
    InMux I__7094 (
            .O(N__34986),
            .I(N__34958));
    InMux I__7093 (
            .O(N__34985),
            .I(N__34958));
    Span4Mux_h I__7092 (
            .O(N__34982),
            .I(N__34955));
    Span4Mux_h I__7091 (
            .O(N__34979),
            .I(N__34950));
    LocalMux I__7090 (
            .O(N__34976),
            .I(N__34950));
    LocalMux I__7089 (
            .O(N__34969),
            .I(N__34945));
    LocalMux I__7088 (
            .O(N__34964),
            .I(N__34942));
    InMux I__7087 (
            .O(N__34963),
            .I(N__34939));
    LocalMux I__7086 (
            .O(N__34958),
            .I(N__34936));
    Span4Mux_v I__7085 (
            .O(N__34955),
            .I(N__34933));
    Span4Mux_v I__7084 (
            .O(N__34950),
            .I(N__34930));
    InMux I__7083 (
            .O(N__34949),
            .I(N__34925));
    InMux I__7082 (
            .O(N__34948),
            .I(N__34925));
    Span12Mux_s11_v I__7081 (
            .O(N__34945),
            .I(N__34922));
    Span4Mux_v I__7080 (
            .O(N__34942),
            .I(N__34915));
    LocalMux I__7079 (
            .O(N__34939),
            .I(N__34915));
    Span4Mux_h I__7078 (
            .O(N__34936),
            .I(N__34915));
    Odrv4 I__7077 (
            .O(N__34933),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7076 (
            .O(N__34930),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    LocalMux I__7075 (
            .O(N__34925),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv12 I__7074 (
            .O(N__34922),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7073 (
            .O(N__34915),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    InMux I__7072 (
            .O(N__34904),
            .I(N__34900));
    InMux I__7071 (
            .O(N__34903),
            .I(N__34897));
    LocalMux I__7070 (
            .O(N__34900),
            .I(N__34894));
    LocalMux I__7069 (
            .O(N__34897),
            .I(N__34888));
    Span4Mux_h I__7068 (
            .O(N__34894),
            .I(N__34888));
    InMux I__7067 (
            .O(N__34893),
            .I(N__34885));
    Span4Mux_v I__7066 (
            .O(N__34888),
            .I(N__34880));
    LocalMux I__7065 (
            .O(N__34885),
            .I(N__34880));
    Odrv4 I__7064 (
            .O(N__34880),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    InMux I__7063 (
            .O(N__34877),
            .I(N__34874));
    LocalMux I__7062 (
            .O(N__34874),
            .I(N__34870));
    InMux I__7061 (
            .O(N__34873),
            .I(N__34867));
    Span4Mux_h I__7060 (
            .O(N__34870),
            .I(N__34864));
    LocalMux I__7059 (
            .O(N__34867),
            .I(N__34861));
    Odrv4 I__7058 (
            .O(N__34864),
            .I(\phase_controller_inst1.stoper_hc.un1_N_4 ));
    Odrv12 I__7057 (
            .O(N__34861),
            .I(\phase_controller_inst1.stoper_hc.un1_N_4 ));
    InMux I__7056 (
            .O(N__34856),
            .I(N__34853));
    LocalMux I__7055 (
            .O(N__34853),
            .I(N__34850));
    Span4Mux_h I__7054 (
            .O(N__34850),
            .I(N__34847));
    Odrv4 I__7053 (
            .O(N__34847),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0 ));
    InMux I__7052 (
            .O(N__34844),
            .I(N__34840));
    InMux I__7051 (
            .O(N__34843),
            .I(N__34837));
    LocalMux I__7050 (
            .O(N__34840),
            .I(N__34834));
    LocalMux I__7049 (
            .O(N__34837),
            .I(N__34831));
    Span4Mux_h I__7048 (
            .O(N__34834),
            .I(N__34828));
    Odrv4 I__7047 (
            .O(N__34831),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7046 (
            .O(N__34828),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__7045 (
            .O(N__34823),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0_cascade_ ));
    CascadeMux I__7044 (
            .O(N__34820),
            .I(N__34817));
    InMux I__7043 (
            .O(N__34817),
            .I(N__34813));
    InMux I__7042 (
            .O(N__34816),
            .I(N__34810));
    LocalMux I__7041 (
            .O(N__34813),
            .I(N__34804));
    LocalMux I__7040 (
            .O(N__34810),
            .I(N__34801));
    InMux I__7039 (
            .O(N__34809),
            .I(N__34796));
    InMux I__7038 (
            .O(N__34808),
            .I(N__34796));
    CascadeMux I__7037 (
            .O(N__34807),
            .I(N__34793));
    Span4Mux_h I__7036 (
            .O(N__34804),
            .I(N__34786));
    Span4Mux_h I__7035 (
            .O(N__34801),
            .I(N__34786));
    LocalMux I__7034 (
            .O(N__34796),
            .I(N__34786));
    InMux I__7033 (
            .O(N__34793),
            .I(N__34783));
    Span4Mux_v I__7032 (
            .O(N__34786),
            .I(N__34780));
    LocalMux I__7031 (
            .O(N__34783),
            .I(measured_delay_hc_16));
    Odrv4 I__7030 (
            .O(N__34780),
            .I(measured_delay_hc_16));
    InMux I__7029 (
            .O(N__34775),
            .I(N__34772));
    LocalMux I__7028 (
            .O(N__34772),
            .I(N__34765));
    InMux I__7027 (
            .O(N__34771),
            .I(N__34758));
    InMux I__7026 (
            .O(N__34770),
            .I(N__34758));
    InMux I__7025 (
            .O(N__34769),
            .I(N__34758));
    InMux I__7024 (
            .O(N__34768),
            .I(N__34755));
    Span4Mux_h I__7023 (
            .O(N__34765),
            .I(N__34752));
    LocalMux I__7022 (
            .O(N__34758),
            .I(N__34749));
    LocalMux I__7021 (
            .O(N__34755),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0 ));
    Odrv4 I__7020 (
            .O(N__34752),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0 ));
    Odrv4 I__7019 (
            .O(N__34749),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0 ));
    CascadeMux I__7018 (
            .O(N__34742),
            .I(N__34738));
    CascadeMux I__7017 (
            .O(N__34741),
            .I(N__34733));
    InMux I__7016 (
            .O(N__34738),
            .I(N__34729));
    InMux I__7015 (
            .O(N__34737),
            .I(N__34726));
    InMux I__7014 (
            .O(N__34736),
            .I(N__34721));
    InMux I__7013 (
            .O(N__34733),
            .I(N__34721));
    CascadeMux I__7012 (
            .O(N__34732),
            .I(N__34718));
    LocalMux I__7011 (
            .O(N__34729),
            .I(N__34715));
    LocalMux I__7010 (
            .O(N__34726),
            .I(N__34712));
    LocalMux I__7009 (
            .O(N__34721),
            .I(N__34709));
    InMux I__7008 (
            .O(N__34718),
            .I(N__34706));
    Span12Mux_v I__7007 (
            .O(N__34715),
            .I(N__34703));
    Span4Mux_v I__7006 (
            .O(N__34712),
            .I(N__34698));
    Span4Mux_h I__7005 (
            .O(N__34709),
            .I(N__34698));
    LocalMux I__7004 (
            .O(N__34706),
            .I(measured_delay_hc_17));
    Odrv12 I__7003 (
            .O(N__34703),
            .I(measured_delay_hc_17));
    Odrv4 I__7002 (
            .O(N__34698),
            .I(measured_delay_hc_17));
    CascadeMux I__7001 (
            .O(N__34691),
            .I(N__34688));
    InMux I__7000 (
            .O(N__34688),
            .I(N__34685));
    LocalMux I__6999 (
            .O(N__34685),
            .I(N__34682));
    Span12Mux_s8_v I__6998 (
            .O(N__34682),
            .I(N__34677));
    InMux I__6997 (
            .O(N__34681),
            .I(N__34674));
    InMux I__6996 (
            .O(N__34680),
            .I(N__34669));
    Span12Mux_h I__6995 (
            .O(N__34677),
            .I(N__34664));
    LocalMux I__6994 (
            .O(N__34674),
            .I(N__34664));
    InMux I__6993 (
            .O(N__34673),
            .I(N__34661));
    InMux I__6992 (
            .O(N__34672),
            .I(N__34658));
    LocalMux I__6991 (
            .O(N__34669),
            .I(measured_delay_hc_10));
    Odrv12 I__6990 (
            .O(N__34664),
            .I(measured_delay_hc_10));
    LocalMux I__6989 (
            .O(N__34661),
            .I(measured_delay_hc_10));
    LocalMux I__6988 (
            .O(N__34658),
            .I(measured_delay_hc_10));
    InMux I__6987 (
            .O(N__34649),
            .I(N__34645));
    InMux I__6986 (
            .O(N__34648),
            .I(N__34642));
    LocalMux I__6985 (
            .O(N__34645),
            .I(N__34637));
    LocalMux I__6984 (
            .O(N__34642),
            .I(N__34633));
    InMux I__6983 (
            .O(N__34641),
            .I(N__34630));
    InMux I__6982 (
            .O(N__34640),
            .I(N__34627));
    Span4Mux_v I__6981 (
            .O(N__34637),
            .I(N__34624));
    InMux I__6980 (
            .O(N__34636),
            .I(N__34621));
    Span4Mux_v I__6979 (
            .O(N__34633),
            .I(N__34616));
    LocalMux I__6978 (
            .O(N__34630),
            .I(N__34616));
    LocalMux I__6977 (
            .O(N__34627),
            .I(measured_delay_hc_11));
    Odrv4 I__6976 (
            .O(N__34624),
            .I(measured_delay_hc_11));
    LocalMux I__6975 (
            .O(N__34621),
            .I(measured_delay_hc_11));
    Odrv4 I__6974 (
            .O(N__34616),
            .I(measured_delay_hc_11));
    CascadeMux I__6973 (
            .O(N__34607),
            .I(N__34603));
    CascadeMux I__6972 (
            .O(N__34606),
            .I(N__34600));
    InMux I__6971 (
            .O(N__34603),
            .I(N__34597));
    InMux I__6970 (
            .O(N__34600),
            .I(N__34592));
    LocalMux I__6969 (
            .O(N__34597),
            .I(N__34589));
    InMux I__6968 (
            .O(N__34596),
            .I(N__34586));
    InMux I__6967 (
            .O(N__34595),
            .I(N__34583));
    LocalMux I__6966 (
            .O(N__34592),
            .I(N__34578));
    Span4Mux_v I__6965 (
            .O(N__34589),
            .I(N__34578));
    LocalMux I__6964 (
            .O(N__34586),
            .I(N__34575));
    LocalMux I__6963 (
            .O(N__34583),
            .I(N__34572));
    Odrv4 I__6962 (
            .O(N__34578),
            .I(measured_delay_hc_2));
    Odrv12 I__6961 (
            .O(N__34575),
            .I(measured_delay_hc_2));
    Odrv4 I__6960 (
            .O(N__34572),
            .I(measured_delay_hc_2));
    CascadeMux I__6959 (
            .O(N__34565),
            .I(N__34562));
    InMux I__6958 (
            .O(N__34562),
            .I(N__34558));
    InMux I__6957 (
            .O(N__34561),
            .I(N__34553));
    LocalMux I__6956 (
            .O(N__34558),
            .I(N__34550));
    InMux I__6955 (
            .O(N__34557),
            .I(N__34547));
    InMux I__6954 (
            .O(N__34556),
            .I(N__34544));
    LocalMux I__6953 (
            .O(N__34553),
            .I(N__34540));
    Span4Mux_v I__6952 (
            .O(N__34550),
            .I(N__34533));
    LocalMux I__6951 (
            .O(N__34547),
            .I(N__34533));
    LocalMux I__6950 (
            .O(N__34544),
            .I(N__34533));
    InMux I__6949 (
            .O(N__34543),
            .I(N__34530));
    Span4Mux_h I__6948 (
            .O(N__34540),
            .I(N__34527));
    Span4Mux_v I__6947 (
            .O(N__34533),
            .I(N__34524));
    LocalMux I__6946 (
            .O(N__34530),
            .I(measured_delay_hc_7));
    Odrv4 I__6945 (
            .O(N__34527),
            .I(measured_delay_hc_7));
    Odrv4 I__6944 (
            .O(N__34524),
            .I(measured_delay_hc_7));
    InMux I__6943 (
            .O(N__34517),
            .I(N__34514));
    LocalMux I__6942 (
            .O(N__34514),
            .I(N__34508));
    InMux I__6941 (
            .O(N__34513),
            .I(N__34505));
    InMux I__6940 (
            .O(N__34512),
            .I(N__34502));
    InMux I__6939 (
            .O(N__34511),
            .I(N__34499));
    Span12Mux_h I__6938 (
            .O(N__34508),
            .I(N__34492));
    LocalMux I__6937 (
            .O(N__34505),
            .I(N__34492));
    LocalMux I__6936 (
            .O(N__34502),
            .I(N__34492));
    LocalMux I__6935 (
            .O(N__34499),
            .I(measured_delay_hc_5));
    Odrv12 I__6934 (
            .O(N__34492),
            .I(measured_delay_hc_5));
    InMux I__6933 (
            .O(N__34487),
            .I(N__34483));
    InMux I__6932 (
            .O(N__34486),
            .I(N__34480));
    LocalMux I__6931 (
            .O(N__34483),
            .I(N__34477));
    LocalMux I__6930 (
            .O(N__34480),
            .I(measured_delay_hc_23));
    Odrv4 I__6929 (
            .O(N__34477),
            .I(measured_delay_hc_23));
    InMux I__6928 (
            .O(N__34472),
            .I(N__34469));
    LocalMux I__6927 (
            .O(N__34469),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3 ));
    CascadeMux I__6926 (
            .O(N__34466),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__6925 (
            .O(N__34463),
            .I(N__34460));
    LocalMux I__6924 (
            .O(N__34460),
            .I(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ));
    InMux I__6923 (
            .O(N__34457),
            .I(N__34454));
    LocalMux I__6922 (
            .O(N__34454),
            .I(N__34447));
    InMux I__6921 (
            .O(N__34453),
            .I(N__34444));
    InMux I__6920 (
            .O(N__34452),
            .I(N__34439));
    InMux I__6919 (
            .O(N__34451),
            .I(N__34439));
    CascadeMux I__6918 (
            .O(N__34450),
            .I(N__34436));
    Span4Mux_v I__6917 (
            .O(N__34447),
            .I(N__34431));
    LocalMux I__6916 (
            .O(N__34444),
            .I(N__34431));
    LocalMux I__6915 (
            .O(N__34439),
            .I(N__34428));
    InMux I__6914 (
            .O(N__34436),
            .I(N__34425));
    Span4Mux_v I__6913 (
            .O(N__34431),
            .I(N__34422));
    Span4Mux_h I__6912 (
            .O(N__34428),
            .I(N__34419));
    LocalMux I__6911 (
            .O(N__34425),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__6910 (
            .O(N__34422),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__6909 (
            .O(N__34419),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    InMux I__6908 (
            .O(N__34412),
            .I(N__34407));
    InMux I__6907 (
            .O(N__34411),
            .I(N__34404));
    InMux I__6906 (
            .O(N__34410),
            .I(N__34401));
    LocalMux I__6905 (
            .O(N__34407),
            .I(N__34396));
    LocalMux I__6904 (
            .O(N__34404),
            .I(N__34396));
    LocalMux I__6903 (
            .O(N__34401),
            .I(N__34393));
    Span4Mux_v I__6902 (
            .O(N__34396),
            .I(N__34390));
    Span12Mux_v I__6901 (
            .O(N__34393),
            .I(N__34387));
    Span4Mux_h I__6900 (
            .O(N__34390),
            .I(N__34384));
    Odrv12 I__6899 (
            .O(N__34387),
            .I(il_max_comp1_D2));
    Odrv4 I__6898 (
            .O(N__34384),
            .I(il_max_comp1_D2));
    InMux I__6897 (
            .O(N__34379),
            .I(N__34375));
    CascadeMux I__6896 (
            .O(N__34378),
            .I(N__34372));
    LocalMux I__6895 (
            .O(N__34375),
            .I(N__34368));
    InMux I__6894 (
            .O(N__34372),
            .I(N__34363));
    InMux I__6893 (
            .O(N__34371),
            .I(N__34363));
    Odrv4 I__6892 (
            .O(N__34368),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6891 (
            .O(N__34363),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__6890 (
            .O(N__34358),
            .I(N__34355));
    InMux I__6889 (
            .O(N__34355),
            .I(N__34352));
    LocalMux I__6888 (
            .O(N__34352),
            .I(N__34349));
    Odrv4 I__6887 (
            .O(N__34349),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__6886 (
            .O(N__34346),
            .I(N__34342));
    InMux I__6885 (
            .O(N__34345),
            .I(N__34337));
    LocalMux I__6884 (
            .O(N__34342),
            .I(N__34334));
    InMux I__6883 (
            .O(N__34341),
            .I(N__34329));
    InMux I__6882 (
            .O(N__34340),
            .I(N__34329));
    LocalMux I__6881 (
            .O(N__34337),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__6880 (
            .O(N__34334),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__6879 (
            .O(N__34329),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__6878 (
            .O(N__34322),
            .I(N__34318));
    InMux I__6877 (
            .O(N__34321),
            .I(N__34315));
    LocalMux I__6876 (
            .O(N__34318),
            .I(N__34309));
    LocalMux I__6875 (
            .O(N__34315),
            .I(N__34309));
    InMux I__6874 (
            .O(N__34314),
            .I(N__34306));
    Span4Mux_h I__6873 (
            .O(N__34309),
            .I(N__34303));
    LocalMux I__6872 (
            .O(N__34306),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__6871 (
            .O(N__34303),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    CascadeMux I__6870 (
            .O(N__34298),
            .I(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ));
    InMux I__6869 (
            .O(N__34295),
            .I(N__34287));
    InMux I__6868 (
            .O(N__34294),
            .I(N__34287));
    InMux I__6867 (
            .O(N__34293),
            .I(N__34280));
    InMux I__6866 (
            .O(N__34292),
            .I(N__34280));
    LocalMux I__6865 (
            .O(N__34287),
            .I(N__34277));
    InMux I__6864 (
            .O(N__34286),
            .I(N__34274));
    InMux I__6863 (
            .O(N__34285),
            .I(N__34271));
    LocalMux I__6862 (
            .O(N__34280),
            .I(N__34268));
    Odrv4 I__6861 (
            .O(N__34277),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6860 (
            .O(N__34274),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6859 (
            .O(N__34271),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__6858 (
            .O(N__34268),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__6857 (
            .O(N__34259),
            .I(N__34256));
    LocalMux I__6856 (
            .O(N__34256),
            .I(N__34253));
    Span4Mux_h I__6855 (
            .O(N__34253),
            .I(N__34249));
    InMux I__6854 (
            .O(N__34252),
            .I(N__34245));
    Span4Mux_v I__6853 (
            .O(N__34249),
            .I(N__34242));
    CascadeMux I__6852 (
            .O(N__34248),
            .I(N__34239));
    LocalMux I__6851 (
            .O(N__34245),
            .I(N__34235));
    Sp12to4 I__6850 (
            .O(N__34242),
            .I(N__34232));
    InMux I__6849 (
            .O(N__34239),
            .I(N__34227));
    InMux I__6848 (
            .O(N__34238),
            .I(N__34227));
    Odrv4 I__6847 (
            .O(N__34235),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv12 I__6846 (
            .O(N__34232),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    LocalMux I__6845 (
            .O(N__34227),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    InMux I__6844 (
            .O(N__34220),
            .I(N__34216));
    InMux I__6843 (
            .O(N__34219),
            .I(N__34213));
    LocalMux I__6842 (
            .O(N__34216),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1 ));
    LocalMux I__6841 (
            .O(N__34213),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1 ));
    InMux I__6840 (
            .O(N__34208),
            .I(N__34205));
    LocalMux I__6839 (
            .O(N__34205),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ));
    InMux I__6838 (
            .O(N__34202),
            .I(N__34196));
    InMux I__6837 (
            .O(N__34201),
            .I(N__34196));
    LocalMux I__6836 (
            .O(N__34196),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2 ));
    InMux I__6835 (
            .O(N__34193),
            .I(N__34190));
    LocalMux I__6834 (
            .O(N__34190),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ));
    InMux I__6833 (
            .O(N__34187),
            .I(N__34184));
    LocalMux I__6832 (
            .O(N__34184),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ));
    CascadeMux I__6831 (
            .O(N__34181),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ));
    InMux I__6830 (
            .O(N__34178),
            .I(N__34173));
    InMux I__6829 (
            .O(N__34177),
            .I(N__34170));
    InMux I__6828 (
            .O(N__34176),
            .I(N__34167));
    LocalMux I__6827 (
            .O(N__34173),
            .I(N__34162));
    LocalMux I__6826 (
            .O(N__34170),
            .I(N__34162));
    LocalMux I__6825 (
            .O(N__34167),
            .I(N__34159));
    Span4Mux_h I__6824 (
            .O(N__34162),
            .I(N__34156));
    Span4Mux_h I__6823 (
            .O(N__34159),
            .I(N__34153));
    Sp12to4 I__6822 (
            .O(N__34156),
            .I(N__34150));
    Sp12to4 I__6821 (
            .O(N__34153),
            .I(N__34145));
    Span12Mux_v I__6820 (
            .O(N__34150),
            .I(N__34145));
    Odrv12 I__6819 (
            .O(N__34145),
            .I(il_min_comp1_D2));
    InMux I__6818 (
            .O(N__34142),
            .I(N__34137));
    InMux I__6817 (
            .O(N__34141),
            .I(N__34133));
    InMux I__6816 (
            .O(N__34140),
            .I(N__34130));
    LocalMux I__6815 (
            .O(N__34137),
            .I(N__34127));
    InMux I__6814 (
            .O(N__34136),
            .I(N__34124));
    LocalMux I__6813 (
            .O(N__34133),
            .I(N__34120));
    LocalMux I__6812 (
            .O(N__34130),
            .I(N__34113));
    Span4Mux_v I__6811 (
            .O(N__34127),
            .I(N__34113));
    LocalMux I__6810 (
            .O(N__34124),
            .I(N__34113));
    CascadeMux I__6809 (
            .O(N__34123),
            .I(N__34110));
    Sp12to4 I__6808 (
            .O(N__34120),
            .I(N__34105));
    Sp12to4 I__6807 (
            .O(N__34113),
            .I(N__34105));
    InMux I__6806 (
            .O(N__34110),
            .I(N__34102));
    Span12Mux_s11_v I__6805 (
            .O(N__34105),
            .I(N__34099));
    LocalMux I__6804 (
            .O(N__34102),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__6803 (
            .O(N__34099),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__6802 (
            .O(N__34094),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__6801 (
            .O(N__34091),
            .I(N__34088));
    LocalMux I__6800 (
            .O(N__34088),
            .I(N__34085));
    Odrv4 I__6799 (
            .O(N__34085),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__6798 (
            .O(N__34082),
            .I(N__34079));
    LocalMux I__6797 (
            .O(N__34079),
            .I(N__34076));
    Odrv4 I__6796 (
            .O(N__34076),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    IoInMux I__6795 (
            .O(N__34073),
            .I(N__34070));
    LocalMux I__6794 (
            .O(N__34070),
            .I(s2_phy_c));
    IoInMux I__6793 (
            .O(N__34067),
            .I(N__34064));
    LocalMux I__6792 (
            .O(N__34064),
            .I(N__34061));
    Span4Mux_s3_v I__6791 (
            .O(N__34061),
            .I(N__34058));
    Odrv4 I__6790 (
            .O(N__34058),
            .I(\delay_measurement_inst.delay_hc_timer.N_335_i ));
    InMux I__6789 (
            .O(N__34055),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__6788 (
            .O(N__34052),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__6787 (
            .O(N__34049),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__6786 (
            .O(N__34046),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__6785 (
            .O(N__34043),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__6784 (
            .O(N__34040),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__6783 (
            .O(N__34037),
            .I(N__34034));
    LocalMux I__6782 (
            .O(N__34034),
            .I(N__34031));
    Odrv4 I__6781 (
            .O(N__34031),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__6780 (
            .O(N__34028),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__6779 (
            .O(N__34025),
            .I(bfn_13_26_0_));
    InMux I__6778 (
            .O(N__34022),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__6777 (
            .O(N__34019),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__6776 (
            .O(N__34016),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__6775 (
            .O(N__34013),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__6774 (
            .O(N__34010),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__6773 (
            .O(N__34007),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__6772 (
            .O(N__34004),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__6771 (
            .O(N__34001),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__6770 (
            .O(N__33998),
            .I(bfn_13_25_0_));
    InMux I__6769 (
            .O(N__33995),
            .I(N__33991));
    InMux I__6768 (
            .O(N__33994),
            .I(N__33988));
    LocalMux I__6767 (
            .O(N__33991),
            .I(N__33984));
    LocalMux I__6766 (
            .O(N__33988),
            .I(N__33981));
    InMux I__6765 (
            .O(N__33987),
            .I(N__33978));
    Span4Mux_v I__6764 (
            .O(N__33984),
            .I(N__33975));
    Span4Mux_h I__6763 (
            .O(N__33981),
            .I(N__33972));
    LocalMux I__6762 (
            .O(N__33978),
            .I(N__33969));
    Span4Mux_v I__6761 (
            .O(N__33975),
            .I(N__33966));
    Span4Mux_v I__6760 (
            .O(N__33972),
            .I(N__33961));
    Span4Mux_v I__6759 (
            .O(N__33969),
            .I(N__33961));
    Span4Mux_v I__6758 (
            .O(N__33966),
            .I(N__33958));
    Span4Mux_v I__6757 (
            .O(N__33961),
            .I(N__33955));
    Odrv4 I__6756 (
            .O(N__33958),
            .I(il_min_comp2_D2));
    Odrv4 I__6755 (
            .O(N__33955),
            .I(il_min_comp2_D2));
    InMux I__6754 (
            .O(N__33950),
            .I(N__33946));
    CascadeMux I__6753 (
            .O(N__33949),
            .I(N__33942));
    LocalMux I__6752 (
            .O(N__33946),
            .I(N__33938));
    InMux I__6751 (
            .O(N__33945),
            .I(N__33935));
    InMux I__6750 (
            .O(N__33942),
            .I(N__33930));
    InMux I__6749 (
            .O(N__33941),
            .I(N__33930));
    Span4Mux_h I__6748 (
            .O(N__33938),
            .I(N__33927));
    LocalMux I__6747 (
            .O(N__33935),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__6746 (
            .O(N__33930),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    Odrv4 I__6745 (
            .O(N__33927),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    CascadeMux I__6744 (
            .O(N__33920),
            .I(N__33917));
    InMux I__6743 (
            .O(N__33917),
            .I(N__33914));
    LocalMux I__6742 (
            .O(N__33914),
            .I(N__33911));
    Odrv4 I__6741 (
            .O(N__33911),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    InMux I__6740 (
            .O(N__33908),
            .I(N__33905));
    LocalMux I__6739 (
            .O(N__33905),
            .I(\phase_controller_slave.state_RNIVDE2Z0Z_0 ));
    IoInMux I__6738 (
            .O(N__33902),
            .I(N__33899));
    LocalMux I__6737 (
            .O(N__33899),
            .I(N__33896));
    IoSpan4Mux I__6736 (
            .O(N__33896),
            .I(N__33892));
    InMux I__6735 (
            .O(N__33895),
            .I(N__33889));
    Span4Mux_s3_v I__6734 (
            .O(N__33892),
            .I(N__33884));
    LocalMux I__6733 (
            .O(N__33889),
            .I(N__33884));
    Span4Mux_v I__6732 (
            .O(N__33884),
            .I(N__33880));
    InMux I__6731 (
            .O(N__33883),
            .I(N__33877));
    Odrv4 I__6730 (
            .O(N__33880),
            .I(s3_phy_c));
    LocalMux I__6729 (
            .O(N__33877),
            .I(s3_phy_c));
    CascadeMux I__6728 (
            .O(N__33872),
            .I(N__33868));
    CascadeMux I__6727 (
            .O(N__33871),
            .I(N__33865));
    InMux I__6726 (
            .O(N__33868),
            .I(N__33861));
    InMux I__6725 (
            .O(N__33865),
            .I(N__33856));
    InMux I__6724 (
            .O(N__33864),
            .I(N__33856));
    LocalMux I__6723 (
            .O(N__33861),
            .I(shift_flag_start));
    LocalMux I__6722 (
            .O(N__33856),
            .I(shift_flag_start));
    InMux I__6721 (
            .O(N__33851),
            .I(N__33848));
    LocalMux I__6720 (
            .O(N__33848),
            .I(N__33845));
    Sp12to4 I__6719 (
            .O(N__33845),
            .I(N__33841));
    InMux I__6718 (
            .O(N__33844),
            .I(N__33838));
    Odrv12 I__6717 (
            .O(N__33841),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    LocalMux I__6716 (
            .O(N__33838),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    CascadeMux I__6715 (
            .O(N__33833),
            .I(N__33830));
    InMux I__6714 (
            .O(N__33830),
            .I(N__33827));
    LocalMux I__6713 (
            .O(N__33827),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__6712 (
            .O(N__33824),
            .I(N__33821));
    LocalMux I__6711 (
            .O(N__33821),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    CascadeMux I__6710 (
            .O(N__33818),
            .I(N__33814));
    InMux I__6709 (
            .O(N__33817),
            .I(N__33806));
    InMux I__6708 (
            .O(N__33814),
            .I(N__33806));
    InMux I__6707 (
            .O(N__33813),
            .I(N__33806));
    LocalMux I__6706 (
            .O(N__33806),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__6705 (
            .O(N__33803),
            .I(N__33797));
    InMux I__6704 (
            .O(N__33802),
            .I(N__33797));
    LocalMux I__6703 (
            .O(N__33797),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CascadeMux I__6702 (
            .O(N__33794),
            .I(N__33791));
    InMux I__6701 (
            .O(N__33791),
            .I(N__33788));
    LocalMux I__6700 (
            .O(N__33788),
            .I(N__33785));
    Span4Mux_h I__6699 (
            .O(N__33785),
            .I(N__33782));
    Odrv4 I__6698 (
            .O(N__33782),
            .I(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ));
    CascadeMux I__6697 (
            .O(N__33779),
            .I(N__33775));
    InMux I__6696 (
            .O(N__33778),
            .I(N__33771));
    InMux I__6695 (
            .O(N__33775),
            .I(N__33766));
    InMux I__6694 (
            .O(N__33774),
            .I(N__33766));
    LocalMux I__6693 (
            .O(N__33771),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__6692 (
            .O(N__33766),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__6691 (
            .O(N__33761),
            .I(N__33755));
    InMux I__6690 (
            .O(N__33760),
            .I(N__33755));
    LocalMux I__6689 (
            .O(N__33755),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    CascadeMux I__6688 (
            .O(N__33752),
            .I(\phase_controller_slave.state_RNIVDE2Z0Z_0_cascade_ ));
    InMux I__6687 (
            .O(N__33749),
            .I(N__33746));
    LocalMux I__6686 (
            .O(N__33746),
            .I(N__33743));
    Span4Mux_h I__6685 (
            .O(N__33743),
            .I(N__33739));
    InMux I__6684 (
            .O(N__33742),
            .I(N__33736));
    Odrv4 I__6683 (
            .O(N__33739),
            .I(state_ns_i_a2_1));
    LocalMux I__6682 (
            .O(N__33736),
            .I(state_ns_i_a2_1));
    InMux I__6681 (
            .O(N__33731),
            .I(N__33726));
    InMux I__6680 (
            .O(N__33730),
            .I(N__33723));
    InMux I__6679 (
            .O(N__33729),
            .I(N__33719));
    LocalMux I__6678 (
            .O(N__33726),
            .I(N__33715));
    LocalMux I__6677 (
            .O(N__33723),
            .I(N__33712));
    CascadeMux I__6676 (
            .O(N__33722),
            .I(N__33709));
    LocalMux I__6675 (
            .O(N__33719),
            .I(N__33706));
    InMux I__6674 (
            .O(N__33718),
            .I(N__33703));
    Span4Mux_v I__6673 (
            .O(N__33715),
            .I(N__33700));
    Span4Mux_h I__6672 (
            .O(N__33712),
            .I(N__33697));
    InMux I__6671 (
            .O(N__33709),
            .I(N__33694));
    Span4Mux_h I__6670 (
            .O(N__33706),
            .I(N__33688));
    LocalMux I__6669 (
            .O(N__33703),
            .I(N__33688));
    Span4Mux_h I__6668 (
            .O(N__33700),
            .I(N__33683));
    Span4Mux_v I__6667 (
            .O(N__33697),
            .I(N__33683));
    LocalMux I__6666 (
            .O(N__33694),
            .I(N__33680));
    InMux I__6665 (
            .O(N__33693),
            .I(N__33677));
    Span4Mux_v I__6664 (
            .O(N__33688),
            .I(N__33674));
    Sp12to4 I__6663 (
            .O(N__33683),
            .I(N__33671));
    Span4Mux_h I__6662 (
            .O(N__33680),
            .I(N__33668));
    LocalMux I__6661 (
            .O(N__33677),
            .I(N__33665));
    Span4Mux_h I__6660 (
            .O(N__33674),
            .I(N__33662));
    Span12Mux_v I__6659 (
            .O(N__33671),
            .I(N__33655));
    Sp12to4 I__6658 (
            .O(N__33668),
            .I(N__33655));
    Sp12to4 I__6657 (
            .O(N__33665),
            .I(N__33655));
    Sp12to4 I__6656 (
            .O(N__33662),
            .I(N__33652));
    Span12Mux_v I__6655 (
            .O(N__33655),
            .I(N__33649));
    Span12Mux_v I__6654 (
            .O(N__33652),
            .I(N__33644));
    Span12Mux_h I__6653 (
            .O(N__33649),
            .I(N__33644));
    Odrv12 I__6652 (
            .O(N__33644),
            .I(start_stop_c));
    IoInMux I__6651 (
            .O(N__33641),
            .I(N__33638));
    LocalMux I__6650 (
            .O(N__33638),
            .I(N__33635));
    Span4Mux_s3_v I__6649 (
            .O(N__33635),
            .I(N__33632));
    Span4Mux_h I__6648 (
            .O(N__33632),
            .I(N__33629));
    Span4Mux_v I__6647 (
            .O(N__33629),
            .I(N__33626));
    Span4Mux_v I__6646 (
            .O(N__33626),
            .I(N__33622));
    InMux I__6645 (
            .O(N__33625),
            .I(N__33619));
    Odrv4 I__6644 (
            .O(N__33622),
            .I(s4_phy_c));
    LocalMux I__6643 (
            .O(N__33619),
            .I(s4_phy_c));
    CascadeMux I__6642 (
            .O(N__33614),
            .I(N__33611));
    InMux I__6641 (
            .O(N__33611),
            .I(N__33608));
    LocalMux I__6640 (
            .O(N__33608),
            .I(N__33605));
    Span4Mux_v I__6639 (
            .O(N__33605),
            .I(N__33602));
    Odrv4 I__6638 (
            .O(N__33602),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__6637 (
            .O(N__33599),
            .I(N__33596));
    InMux I__6636 (
            .O(N__33596),
            .I(N__33593));
    LocalMux I__6635 (
            .O(N__33593),
            .I(N__33590));
    Odrv4 I__6634 (
            .O(N__33590),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__6633 (
            .O(N__33587),
            .I(N__33584));
    InMux I__6632 (
            .O(N__33584),
            .I(N__33581));
    LocalMux I__6631 (
            .O(N__33581),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__6630 (
            .O(N__33578),
            .I(N__33575));
    InMux I__6629 (
            .O(N__33575),
            .I(N__33572));
    LocalMux I__6628 (
            .O(N__33572),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CEMux I__6627 (
            .O(N__33569),
            .I(N__33566));
    LocalMux I__6626 (
            .O(N__33566),
            .I(N__33562));
    CEMux I__6625 (
            .O(N__33565),
            .I(N__33558));
    Span4Mux_h I__6624 (
            .O(N__33562),
            .I(N__33553));
    CEMux I__6623 (
            .O(N__33561),
            .I(N__33550));
    LocalMux I__6622 (
            .O(N__33558),
            .I(N__33547));
    CEMux I__6621 (
            .O(N__33557),
            .I(N__33544));
    CEMux I__6620 (
            .O(N__33556),
            .I(N__33541));
    Span4Mux_h I__6619 (
            .O(N__33553),
            .I(N__33537));
    LocalMux I__6618 (
            .O(N__33550),
            .I(N__33534));
    Span4Mux_v I__6617 (
            .O(N__33547),
            .I(N__33529));
    LocalMux I__6616 (
            .O(N__33544),
            .I(N__33529));
    LocalMux I__6615 (
            .O(N__33541),
            .I(N__33526));
    CEMux I__6614 (
            .O(N__33540),
            .I(N__33523));
    Span4Mux_h I__6613 (
            .O(N__33537),
            .I(N__33518));
    Span4Mux_v I__6612 (
            .O(N__33534),
            .I(N__33518));
    Span4Mux_h I__6611 (
            .O(N__33529),
            .I(N__33515));
    Span4Mux_h I__6610 (
            .O(N__33526),
            .I(N__33512));
    LocalMux I__6609 (
            .O(N__33523),
            .I(N__33509));
    Span4Mux_v I__6608 (
            .O(N__33518),
            .I(N__33504));
    Span4Mux_v I__6607 (
            .O(N__33515),
            .I(N__33504));
    Span4Mux_v I__6606 (
            .O(N__33512),
            .I(N__33499));
    Span4Mux_h I__6605 (
            .O(N__33509),
            .I(N__33499));
    Odrv4 I__6604 (
            .O(N__33504),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__6603 (
            .O(N__33499),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__6602 (
            .O(N__33494),
            .I(N__33491));
    InMux I__6601 (
            .O(N__33491),
            .I(N__33488));
    LocalMux I__6600 (
            .O(N__33488),
            .I(N__33485));
    Odrv4 I__6599 (
            .O(N__33485),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__6598 (
            .O(N__33482),
            .I(N__33479));
    LocalMux I__6597 (
            .O(N__33479),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__6596 (
            .O(N__33476),
            .I(N__33473));
    LocalMux I__6595 (
            .O(N__33473),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__6594 (
            .O(N__33470),
            .I(N__33467));
    LocalMux I__6593 (
            .O(N__33467),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__6592 (
            .O(N__33464),
            .I(N__33461));
    InMux I__6591 (
            .O(N__33461),
            .I(N__33458));
    LocalMux I__6590 (
            .O(N__33458),
            .I(N__33455));
    Span4Mux_h I__6589 (
            .O(N__33455),
            .I(N__33452));
    Odrv4 I__6588 (
            .O(N__33452),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__6587 (
            .O(N__33449),
            .I(N__33446));
    LocalMux I__6586 (
            .O(N__33446),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__6585 (
            .O(N__33443),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__6584 (
            .O(N__33440),
            .I(N__33437));
    LocalMux I__6583 (
            .O(N__33437),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__6582 (
            .O(N__33434),
            .I(N__33431));
    InMux I__6581 (
            .O(N__33431),
            .I(N__33428));
    LocalMux I__6580 (
            .O(N__33428),
            .I(N__33425));
    Odrv4 I__6579 (
            .O(N__33425),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__6578 (
            .O(N__33422),
            .I(N__33419));
    LocalMux I__6577 (
            .O(N__33419),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__6576 (
            .O(N__33416),
            .I(N__33413));
    InMux I__6575 (
            .O(N__33413),
            .I(N__33410));
    LocalMux I__6574 (
            .O(N__33410),
            .I(N__33407));
    Span4Mux_v I__6573 (
            .O(N__33407),
            .I(N__33404));
    Span4Mux_v I__6572 (
            .O(N__33404),
            .I(N__33401));
    Span4Mux_h I__6571 (
            .O(N__33401),
            .I(N__33398));
    Span4Mux_h I__6570 (
            .O(N__33398),
            .I(N__33395));
    Odrv4 I__6569 (
            .O(N__33395),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__6568 (
            .O(N__33392),
            .I(N__33389));
    LocalMux I__6567 (
            .O(N__33389),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__6566 (
            .O(N__33386),
            .I(N__33383));
    InMux I__6565 (
            .O(N__33383),
            .I(N__33380));
    LocalMux I__6564 (
            .O(N__33380),
            .I(N__33377));
    Sp12to4 I__6563 (
            .O(N__33377),
            .I(N__33374));
    Span12Mux_h I__6562 (
            .O(N__33374),
            .I(N__33371));
    Odrv12 I__6561 (
            .O(N__33371),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__6560 (
            .O(N__33368),
            .I(N__33365));
    LocalMux I__6559 (
            .O(N__33365),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__6558 (
            .O(N__33362),
            .I(N__33359));
    InMux I__6557 (
            .O(N__33359),
            .I(N__33356));
    LocalMux I__6556 (
            .O(N__33356),
            .I(N__33353));
    Odrv4 I__6555 (
            .O(N__33353),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__6554 (
            .O(N__33350),
            .I(N__33347));
    LocalMux I__6553 (
            .O(N__33347),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__6552 (
            .O(N__33344),
            .I(N__33341));
    LocalMux I__6551 (
            .O(N__33341),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__6550 (
            .O(N__33338),
            .I(N__33335));
    InMux I__6549 (
            .O(N__33335),
            .I(N__33332));
    LocalMux I__6548 (
            .O(N__33332),
            .I(N__33329));
    Span4Mux_v I__6547 (
            .O(N__33329),
            .I(N__33326));
    Odrv4 I__6546 (
            .O(N__33326),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__6545 (
            .O(N__33323),
            .I(N__33320));
    LocalMux I__6544 (
            .O(N__33320),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__6543 (
            .O(N__33317),
            .I(N__33314));
    InMux I__6542 (
            .O(N__33314),
            .I(N__33311));
    LocalMux I__6541 (
            .O(N__33311),
            .I(N__33308));
    Odrv12 I__6540 (
            .O(N__33308),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__6539 (
            .O(N__33305),
            .I(N__33302));
    LocalMux I__6538 (
            .O(N__33302),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__6537 (
            .O(N__33299),
            .I(N__33296));
    LocalMux I__6536 (
            .O(N__33296),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__6535 (
            .O(N__33293),
            .I(N__33290));
    LocalMux I__6534 (
            .O(N__33290),
            .I(N__33287));
    Span4Mux_v I__6533 (
            .O(N__33287),
            .I(N__33284));
    Span4Mux_v I__6532 (
            .O(N__33284),
            .I(N__33281));
    Sp12to4 I__6531 (
            .O(N__33281),
            .I(N__33278));
    Odrv12 I__6530 (
            .O(N__33278),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__6529 (
            .O(N__33275),
            .I(N__33272));
    InMux I__6528 (
            .O(N__33272),
            .I(N__33269));
    LocalMux I__6527 (
            .O(N__33269),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__6526 (
            .O(N__33266),
            .I(N__33263));
    LocalMux I__6525 (
            .O(N__33263),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__6524 (
            .O(N__33260),
            .I(N__33257));
    InMux I__6523 (
            .O(N__33257),
            .I(N__33254));
    LocalMux I__6522 (
            .O(N__33254),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__6521 (
            .O(N__33251),
            .I(N__33248));
    LocalMux I__6520 (
            .O(N__33248),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__6519 (
            .O(N__33245),
            .I(N__33242));
    InMux I__6518 (
            .O(N__33242),
            .I(N__33239));
    LocalMux I__6517 (
            .O(N__33239),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__6516 (
            .O(N__33236),
            .I(N__33233));
    LocalMux I__6515 (
            .O(N__33233),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__6514 (
            .O(N__33230),
            .I(N__33227));
    LocalMux I__6513 (
            .O(N__33227),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__6512 (
            .O(N__33224),
            .I(N__33221));
    InMux I__6511 (
            .O(N__33221),
            .I(N__33218));
    LocalMux I__6510 (
            .O(N__33218),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__6509 (
            .O(N__33215),
            .I(N__33212));
    InMux I__6508 (
            .O(N__33212),
            .I(N__33209));
    LocalMux I__6507 (
            .O(N__33209),
            .I(N__33206));
    Span4Mux_h I__6506 (
            .O(N__33206),
            .I(N__33203));
    Odrv4 I__6505 (
            .O(N__33203),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__6504 (
            .O(N__33200),
            .I(N__33197));
    LocalMux I__6503 (
            .O(N__33197),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__6502 (
            .O(N__33194),
            .I(N__33191));
    InMux I__6501 (
            .O(N__33191),
            .I(N__33188));
    LocalMux I__6500 (
            .O(N__33188),
            .I(N__33185));
    Span4Mux_h I__6499 (
            .O(N__33185),
            .I(N__33182));
    Odrv4 I__6498 (
            .O(N__33182),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    InMux I__6497 (
            .O(N__33179),
            .I(N__33176));
    LocalMux I__6496 (
            .O(N__33176),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__6495 (
            .O(N__33173),
            .I(N__33170));
    InMux I__6494 (
            .O(N__33170),
            .I(N__33167));
    LocalMux I__6493 (
            .O(N__33167),
            .I(N__33164));
    Odrv4 I__6492 (
            .O(N__33164),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__6491 (
            .O(N__33161),
            .I(N__33158));
    LocalMux I__6490 (
            .O(N__33158),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__6489 (
            .O(N__33155),
            .I(N__33152));
    LocalMux I__6488 (
            .O(N__33152),
            .I(N__33149));
    Odrv4 I__6487 (
            .O(N__33149),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ));
    InMux I__6486 (
            .O(N__33146),
            .I(N__33143));
    LocalMux I__6485 (
            .O(N__33143),
            .I(N__33139));
    InMux I__6484 (
            .O(N__33142),
            .I(N__33136));
    Span4Mux_h I__6483 (
            .O(N__33139),
            .I(N__33131));
    LocalMux I__6482 (
            .O(N__33136),
            .I(N__33131));
    Span4Mux_v I__6481 (
            .O(N__33131),
            .I(N__33127));
    InMux I__6480 (
            .O(N__33130),
            .I(N__33124));
    Odrv4 I__6479 (
            .O(N__33127),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ));
    LocalMux I__6478 (
            .O(N__33124),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ));
    InMux I__6477 (
            .O(N__33119),
            .I(N__33116));
    LocalMux I__6476 (
            .O(N__33116),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ));
    InMux I__6475 (
            .O(N__33113),
            .I(N__33110));
    LocalMux I__6474 (
            .O(N__33110),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0 ));
    InMux I__6473 (
            .O(N__33107),
            .I(N__33104));
    LocalMux I__6472 (
            .O(N__33104),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12 ));
    CascadeMux I__6471 (
            .O(N__33101),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_ ));
    CascadeMux I__6470 (
            .O(N__33098),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31_cascade_ ));
    InMux I__6469 (
            .O(N__33095),
            .I(N__33092));
    LocalMux I__6468 (
            .O(N__33092),
            .I(N__33089));
    Span4Mux_h I__6467 (
            .O(N__33089),
            .I(N__33086));
    Odrv4 I__6466 (
            .O(N__33086),
            .I(il_max_comp2_D1));
    InMux I__6465 (
            .O(N__33083),
            .I(N__33070));
    InMux I__6464 (
            .O(N__33082),
            .I(N__33045));
    InMux I__6463 (
            .O(N__33081),
            .I(N__33045));
    InMux I__6462 (
            .O(N__33080),
            .I(N__33045));
    InMux I__6461 (
            .O(N__33079),
            .I(N__33045));
    InMux I__6460 (
            .O(N__33078),
            .I(N__33045));
    InMux I__6459 (
            .O(N__33077),
            .I(N__33045));
    InMux I__6458 (
            .O(N__33076),
            .I(N__33045));
    InMux I__6457 (
            .O(N__33075),
            .I(N__33045));
    InMux I__6456 (
            .O(N__33074),
            .I(N__33042));
    CascadeMux I__6455 (
            .O(N__33073),
            .I(N__33038));
    LocalMux I__6454 (
            .O(N__33070),
            .I(N__33031));
    InMux I__6453 (
            .O(N__33069),
            .I(N__33028));
    InMux I__6452 (
            .O(N__33068),
            .I(N__33015));
    InMux I__6451 (
            .O(N__33067),
            .I(N__33015));
    InMux I__6450 (
            .O(N__33066),
            .I(N__33015));
    InMux I__6449 (
            .O(N__33065),
            .I(N__33015));
    InMux I__6448 (
            .O(N__33064),
            .I(N__33015));
    InMux I__6447 (
            .O(N__33063),
            .I(N__33015));
    InMux I__6446 (
            .O(N__33062),
            .I(N__33012));
    LocalMux I__6445 (
            .O(N__33045),
            .I(N__33000));
    LocalMux I__6444 (
            .O(N__33042),
            .I(N__32997));
    InMux I__6443 (
            .O(N__33041),
            .I(N__32994));
    InMux I__6442 (
            .O(N__33038),
            .I(N__32991));
    InMux I__6441 (
            .O(N__33037),
            .I(N__32982));
    InMux I__6440 (
            .O(N__33036),
            .I(N__32982));
    InMux I__6439 (
            .O(N__33035),
            .I(N__32982));
    InMux I__6438 (
            .O(N__33034),
            .I(N__32982));
    Span4Mux_v I__6437 (
            .O(N__33031),
            .I(N__32979));
    LocalMux I__6436 (
            .O(N__33028),
            .I(N__32976));
    LocalMux I__6435 (
            .O(N__33015),
            .I(N__32971));
    LocalMux I__6434 (
            .O(N__33012),
            .I(N__32971));
    InMux I__6433 (
            .O(N__33011),
            .I(N__32968));
    InMux I__6432 (
            .O(N__33010),
            .I(N__32963));
    InMux I__6431 (
            .O(N__33009),
            .I(N__32963));
    InMux I__6430 (
            .O(N__33008),
            .I(N__32958));
    InMux I__6429 (
            .O(N__33007),
            .I(N__32958));
    InMux I__6428 (
            .O(N__33006),
            .I(N__32955));
    InMux I__6427 (
            .O(N__33005),
            .I(N__32950));
    InMux I__6426 (
            .O(N__33004),
            .I(N__32950));
    InMux I__6425 (
            .O(N__33003),
            .I(N__32947));
    Span4Mux_h I__6424 (
            .O(N__33000),
            .I(N__32944));
    Span4Mux_h I__6423 (
            .O(N__32997),
            .I(N__32939));
    LocalMux I__6422 (
            .O(N__32994),
            .I(N__32939));
    LocalMux I__6421 (
            .O(N__32991),
            .I(N__32926));
    LocalMux I__6420 (
            .O(N__32982),
            .I(N__32926));
    Span4Mux_h I__6419 (
            .O(N__32979),
            .I(N__32926));
    Span4Mux_v I__6418 (
            .O(N__32976),
            .I(N__32926));
    Span4Mux_v I__6417 (
            .O(N__32971),
            .I(N__32926));
    LocalMux I__6416 (
            .O(N__32968),
            .I(N__32926));
    LocalMux I__6415 (
            .O(N__32963),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6414 (
            .O(N__32958),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6413 (
            .O(N__32955),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6412 (
            .O(N__32950),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6411 (
            .O(N__32947),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__6410 (
            .O(N__32944),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__6409 (
            .O(N__32939),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__6408 (
            .O(N__32926),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__6407 (
            .O(N__32909),
            .I(N__32904));
    InMux I__6406 (
            .O(N__32908),
            .I(N__32901));
    CascadeMux I__6405 (
            .O(N__32907),
            .I(N__32892));
    LocalMux I__6404 (
            .O(N__32904),
            .I(N__32888));
    LocalMux I__6403 (
            .O(N__32901),
            .I(N__32885));
    InMux I__6402 (
            .O(N__32900),
            .I(N__32882));
    InMux I__6401 (
            .O(N__32899),
            .I(N__32870));
    InMux I__6400 (
            .O(N__32898),
            .I(N__32870));
    InMux I__6399 (
            .O(N__32897),
            .I(N__32870));
    InMux I__6398 (
            .O(N__32896),
            .I(N__32870));
    InMux I__6397 (
            .O(N__32895),
            .I(N__32870));
    InMux I__6396 (
            .O(N__32892),
            .I(N__32865));
    InMux I__6395 (
            .O(N__32891),
            .I(N__32865));
    Span4Mux_v I__6394 (
            .O(N__32888),
            .I(N__32852));
    Span4Mux_h I__6393 (
            .O(N__32885),
            .I(N__32852));
    LocalMux I__6392 (
            .O(N__32882),
            .I(N__32852));
    InMux I__6391 (
            .O(N__32881),
            .I(N__32849));
    LocalMux I__6390 (
            .O(N__32870),
            .I(N__32846));
    LocalMux I__6389 (
            .O(N__32865),
            .I(N__32843));
    CascadeMux I__6388 (
            .O(N__32864),
            .I(N__32831));
    CascadeMux I__6387 (
            .O(N__32863),
            .I(N__32827));
    CascadeMux I__6386 (
            .O(N__32862),
            .I(N__32822));
    CascadeMux I__6385 (
            .O(N__32861),
            .I(N__32819));
    CascadeMux I__6384 (
            .O(N__32860),
            .I(N__32816));
    CascadeMux I__6383 (
            .O(N__32859),
            .I(N__32812));
    Span4Mux_h I__6382 (
            .O(N__32852),
            .I(N__32807));
    LocalMux I__6381 (
            .O(N__32849),
            .I(N__32804));
    Span4Mux_v I__6380 (
            .O(N__32846),
            .I(N__32799));
    Span4Mux_h I__6379 (
            .O(N__32843),
            .I(N__32799));
    InMux I__6378 (
            .O(N__32842),
            .I(N__32790));
    InMux I__6377 (
            .O(N__32841),
            .I(N__32790));
    InMux I__6376 (
            .O(N__32840),
            .I(N__32790));
    InMux I__6375 (
            .O(N__32839),
            .I(N__32790));
    InMux I__6374 (
            .O(N__32838),
            .I(N__32783));
    InMux I__6373 (
            .O(N__32837),
            .I(N__32783));
    InMux I__6372 (
            .O(N__32836),
            .I(N__32783));
    InMux I__6371 (
            .O(N__32835),
            .I(N__32770));
    InMux I__6370 (
            .O(N__32834),
            .I(N__32770));
    InMux I__6369 (
            .O(N__32831),
            .I(N__32770));
    InMux I__6368 (
            .O(N__32830),
            .I(N__32770));
    InMux I__6367 (
            .O(N__32827),
            .I(N__32770));
    InMux I__6366 (
            .O(N__32826),
            .I(N__32770));
    InMux I__6365 (
            .O(N__32825),
            .I(N__32753));
    InMux I__6364 (
            .O(N__32822),
            .I(N__32753));
    InMux I__6363 (
            .O(N__32819),
            .I(N__32753));
    InMux I__6362 (
            .O(N__32816),
            .I(N__32753));
    InMux I__6361 (
            .O(N__32815),
            .I(N__32753));
    InMux I__6360 (
            .O(N__32812),
            .I(N__32753));
    InMux I__6359 (
            .O(N__32811),
            .I(N__32753));
    InMux I__6358 (
            .O(N__32810),
            .I(N__32753));
    Odrv4 I__6357 (
            .O(N__32807),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__6356 (
            .O(N__32804),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__6355 (
            .O(N__32799),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__6354 (
            .O(N__32790),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__6353 (
            .O(N__32783),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__6352 (
            .O(N__32770),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__6351 (
            .O(N__32753),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    CascadeMux I__6350 (
            .O(N__32738),
            .I(N__32735));
    InMux I__6349 (
            .O(N__32735),
            .I(N__32732));
    LocalMux I__6348 (
            .O(N__32732),
            .I(N__32729));
    Span4Mux_h I__6347 (
            .O(N__32729),
            .I(N__32726));
    Odrv4 I__6346 (
            .O(N__32726),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__6345 (
            .O(N__32723),
            .I(N__32717));
    InMux I__6344 (
            .O(N__32722),
            .I(N__32698));
    InMux I__6343 (
            .O(N__32721),
            .I(N__32698));
    InMux I__6342 (
            .O(N__32720),
            .I(N__32695));
    LocalMux I__6341 (
            .O(N__32717),
            .I(N__32688));
    InMux I__6340 (
            .O(N__32716),
            .I(N__32671));
    InMux I__6339 (
            .O(N__32715),
            .I(N__32671));
    InMux I__6338 (
            .O(N__32714),
            .I(N__32671));
    InMux I__6337 (
            .O(N__32713),
            .I(N__32671));
    InMux I__6336 (
            .O(N__32712),
            .I(N__32671));
    InMux I__6335 (
            .O(N__32711),
            .I(N__32671));
    InMux I__6334 (
            .O(N__32710),
            .I(N__32671));
    InMux I__6333 (
            .O(N__32709),
            .I(N__32671));
    InMux I__6332 (
            .O(N__32708),
            .I(N__32658));
    InMux I__6331 (
            .O(N__32707),
            .I(N__32658));
    InMux I__6330 (
            .O(N__32706),
            .I(N__32658));
    InMux I__6329 (
            .O(N__32705),
            .I(N__32658));
    InMux I__6328 (
            .O(N__32704),
            .I(N__32658));
    InMux I__6327 (
            .O(N__32703),
            .I(N__32658));
    LocalMux I__6326 (
            .O(N__32698),
            .I(N__32648));
    LocalMux I__6325 (
            .O(N__32695),
            .I(N__32648));
    InMux I__6324 (
            .O(N__32694),
            .I(N__32639));
    InMux I__6323 (
            .O(N__32693),
            .I(N__32639));
    InMux I__6322 (
            .O(N__32692),
            .I(N__32639));
    InMux I__6321 (
            .O(N__32691),
            .I(N__32639));
    Span4Mux_h I__6320 (
            .O(N__32688),
            .I(N__32635));
    LocalMux I__6319 (
            .O(N__32671),
            .I(N__32632));
    LocalMux I__6318 (
            .O(N__32658),
            .I(N__32629));
    InMux I__6317 (
            .O(N__32657),
            .I(N__32618));
    InMux I__6316 (
            .O(N__32656),
            .I(N__32618));
    InMux I__6315 (
            .O(N__32655),
            .I(N__32618));
    InMux I__6314 (
            .O(N__32654),
            .I(N__32618));
    InMux I__6313 (
            .O(N__32653),
            .I(N__32618));
    Span4Mux_v I__6312 (
            .O(N__32648),
            .I(N__32613));
    LocalMux I__6311 (
            .O(N__32639),
            .I(N__32613));
    InMux I__6310 (
            .O(N__32638),
            .I(N__32610));
    Odrv4 I__6309 (
            .O(N__32635),
            .I(\current_shift_inst.PI_CTRL.N_79 ));
    Odrv4 I__6308 (
            .O(N__32632),
            .I(\current_shift_inst.PI_CTRL.N_79 ));
    Odrv4 I__6307 (
            .O(N__32629),
            .I(\current_shift_inst.PI_CTRL.N_79 ));
    LocalMux I__6306 (
            .O(N__32618),
            .I(\current_shift_inst.PI_CTRL.N_79 ));
    Odrv4 I__6305 (
            .O(N__32613),
            .I(\current_shift_inst.PI_CTRL.N_79 ));
    LocalMux I__6304 (
            .O(N__32610),
            .I(\current_shift_inst.PI_CTRL.N_79 ));
    InMux I__6303 (
            .O(N__32597),
            .I(N__32593));
    InMux I__6302 (
            .O(N__32596),
            .I(N__32590));
    LocalMux I__6301 (
            .O(N__32593),
            .I(N__32585));
    LocalMux I__6300 (
            .O(N__32590),
            .I(N__32582));
    InMux I__6299 (
            .O(N__32589),
            .I(N__32579));
    InMux I__6298 (
            .O(N__32588),
            .I(N__32576));
    Span4Mux_h I__6297 (
            .O(N__32585),
            .I(N__32573));
    Span12Mux_v I__6296 (
            .O(N__32582),
            .I(N__32566));
    LocalMux I__6295 (
            .O(N__32579),
            .I(N__32566));
    LocalMux I__6294 (
            .O(N__32576),
            .I(N__32566));
    Odrv4 I__6293 (
            .O(N__32573),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__6292 (
            .O(N__32566),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    CEMux I__6291 (
            .O(N__32561),
            .I(N__32556));
    CEMux I__6290 (
            .O(N__32560),
            .I(N__32544));
    CEMux I__6289 (
            .O(N__32559),
            .I(N__32541));
    LocalMux I__6288 (
            .O(N__32556),
            .I(N__32537));
    CEMux I__6287 (
            .O(N__32555),
            .I(N__32534));
    CEMux I__6286 (
            .O(N__32554),
            .I(N__32531));
    CEMux I__6285 (
            .O(N__32553),
            .I(N__32527));
    CEMux I__6284 (
            .O(N__32552),
            .I(N__32524));
    CEMux I__6283 (
            .O(N__32551),
            .I(N__32521));
    CEMux I__6282 (
            .O(N__32550),
            .I(N__32518));
    CEMux I__6281 (
            .O(N__32549),
            .I(N__32515));
    CEMux I__6280 (
            .O(N__32548),
            .I(N__32510));
    CEMux I__6279 (
            .O(N__32547),
            .I(N__32507));
    LocalMux I__6278 (
            .O(N__32544),
            .I(N__32504));
    LocalMux I__6277 (
            .O(N__32541),
            .I(N__32501));
    CEMux I__6276 (
            .O(N__32540),
            .I(N__32498));
    Span4Mux_h I__6275 (
            .O(N__32537),
            .I(N__32492));
    LocalMux I__6274 (
            .O(N__32534),
            .I(N__32492));
    LocalMux I__6273 (
            .O(N__32531),
            .I(N__32486));
    CEMux I__6272 (
            .O(N__32530),
            .I(N__32481));
    LocalMux I__6271 (
            .O(N__32527),
            .I(N__32477));
    LocalMux I__6270 (
            .O(N__32524),
            .I(N__32470));
    LocalMux I__6269 (
            .O(N__32521),
            .I(N__32470));
    LocalMux I__6268 (
            .O(N__32518),
            .I(N__32470));
    LocalMux I__6267 (
            .O(N__32515),
            .I(N__32467));
    CEMux I__6266 (
            .O(N__32514),
            .I(N__32464));
    CEMux I__6265 (
            .O(N__32513),
            .I(N__32461));
    LocalMux I__6264 (
            .O(N__32510),
            .I(N__32456));
    LocalMux I__6263 (
            .O(N__32507),
            .I(N__32456));
    Span4Mux_v I__6262 (
            .O(N__32504),
            .I(N__32453));
    Span4Mux_v I__6261 (
            .O(N__32501),
            .I(N__32448));
    LocalMux I__6260 (
            .O(N__32498),
            .I(N__32448));
    CEMux I__6259 (
            .O(N__32497),
            .I(N__32445));
    Span4Mux_h I__6258 (
            .O(N__32492),
            .I(N__32442));
    CEMux I__6257 (
            .O(N__32491),
            .I(N__32439));
    CEMux I__6256 (
            .O(N__32490),
            .I(N__32436));
    CEMux I__6255 (
            .O(N__32489),
            .I(N__32433));
    Span4Mux_h I__6254 (
            .O(N__32486),
            .I(N__32429));
    CEMux I__6253 (
            .O(N__32485),
            .I(N__32426));
    CEMux I__6252 (
            .O(N__32484),
            .I(N__32423));
    LocalMux I__6251 (
            .O(N__32481),
            .I(N__32420));
    CEMux I__6250 (
            .O(N__32480),
            .I(N__32417));
    Span4Mux_v I__6249 (
            .O(N__32477),
            .I(N__32414));
    Span4Mux_v I__6248 (
            .O(N__32470),
            .I(N__32411));
    Span4Mux_h I__6247 (
            .O(N__32467),
            .I(N__32404));
    LocalMux I__6246 (
            .O(N__32464),
            .I(N__32404));
    LocalMux I__6245 (
            .O(N__32461),
            .I(N__32404));
    Span4Mux_v I__6244 (
            .O(N__32456),
            .I(N__32401));
    Span4Mux_h I__6243 (
            .O(N__32453),
            .I(N__32396));
    Span4Mux_h I__6242 (
            .O(N__32448),
            .I(N__32396));
    LocalMux I__6241 (
            .O(N__32445),
            .I(N__32393));
    Span4Mux_h I__6240 (
            .O(N__32442),
            .I(N__32384));
    LocalMux I__6239 (
            .O(N__32439),
            .I(N__32384));
    LocalMux I__6238 (
            .O(N__32436),
            .I(N__32384));
    LocalMux I__6237 (
            .O(N__32433),
            .I(N__32384));
    CEMux I__6236 (
            .O(N__32432),
            .I(N__32381));
    Span4Mux_h I__6235 (
            .O(N__32429),
            .I(N__32376));
    LocalMux I__6234 (
            .O(N__32426),
            .I(N__32376));
    LocalMux I__6233 (
            .O(N__32423),
            .I(N__32373));
    Span12Mux_v I__6232 (
            .O(N__32420),
            .I(N__32370));
    LocalMux I__6231 (
            .O(N__32417),
            .I(N__32367));
    Span4Mux_h I__6230 (
            .O(N__32414),
            .I(N__32358));
    Span4Mux_h I__6229 (
            .O(N__32411),
            .I(N__32358));
    Span4Mux_v I__6228 (
            .O(N__32404),
            .I(N__32358));
    Span4Mux_s3_h I__6227 (
            .O(N__32401),
            .I(N__32358));
    Span4Mux_h I__6226 (
            .O(N__32396),
            .I(N__32349));
    Span4Mux_v I__6225 (
            .O(N__32393),
            .I(N__32349));
    Span4Mux_v I__6224 (
            .O(N__32384),
            .I(N__32349));
    LocalMux I__6223 (
            .O(N__32381),
            .I(N__32349));
    Span4Mux_h I__6222 (
            .O(N__32376),
            .I(N__32344));
    Span4Mux_h I__6221 (
            .O(N__32373),
            .I(N__32344));
    Odrv12 I__6220 (
            .O(N__32370),
            .I(N_605_g));
    Odrv12 I__6219 (
            .O(N__32367),
            .I(N_605_g));
    Odrv4 I__6218 (
            .O(N__32358),
            .I(N_605_g));
    Odrv4 I__6217 (
            .O(N__32349),
            .I(N_605_g));
    Odrv4 I__6216 (
            .O(N__32344),
            .I(N_605_g));
    InMux I__6215 (
            .O(N__32333),
            .I(N__32330));
    LocalMux I__6214 (
            .O(N__32330),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1 ));
    IoInMux I__6213 (
            .O(N__32327),
            .I(N__32324));
    LocalMux I__6212 (
            .O(N__32324),
            .I(N__32321));
    Span4Mux_s3_v I__6211 (
            .O(N__32321),
            .I(N__32318));
    Span4Mux_h I__6210 (
            .O(N__32318),
            .I(N__32314));
    InMux I__6209 (
            .O(N__32317),
            .I(N__32311));
    Odrv4 I__6208 (
            .O(N__32314),
            .I(s1_phy_c));
    LocalMux I__6207 (
            .O(N__32311),
            .I(s1_phy_c));
    CascadeMux I__6206 (
            .O(N__32306),
            .I(N__32302));
    CascadeMux I__6205 (
            .O(N__32305),
            .I(N__32299));
    InMux I__6204 (
            .O(N__32302),
            .I(N__32296));
    InMux I__6203 (
            .O(N__32299),
            .I(N__32293));
    LocalMux I__6202 (
            .O(N__32296),
            .I(N__32289));
    LocalMux I__6201 (
            .O(N__32293),
            .I(N__32286));
    CascadeMux I__6200 (
            .O(N__32292),
            .I(N__32283));
    Span4Mux_v I__6199 (
            .O(N__32289),
            .I(N__32280));
    Span4Mux_v I__6198 (
            .O(N__32286),
            .I(N__32277));
    InMux I__6197 (
            .O(N__32283),
            .I(N__32274));
    Odrv4 I__6196 (
            .O(N__32280),
            .I(\current_shift_inst.S3_riseZ0 ));
    Odrv4 I__6195 (
            .O(N__32277),
            .I(\current_shift_inst.S3_riseZ0 ));
    LocalMux I__6194 (
            .O(N__32274),
            .I(\current_shift_inst.S3_riseZ0 ));
    InMux I__6193 (
            .O(N__32267),
            .I(N__32264));
    LocalMux I__6192 (
            .O(N__32264),
            .I(\current_shift_inst.S3_sync_prevZ0 ));
    InMux I__6191 (
            .O(N__32261),
            .I(N__32258));
    LocalMux I__6190 (
            .O(N__32258),
            .I(\current_shift_inst.S3_syncZ0Z0 ));
    InMux I__6189 (
            .O(N__32255),
            .I(N__32249));
    InMux I__6188 (
            .O(N__32254),
            .I(N__32249));
    LocalMux I__6187 (
            .O(N__32249),
            .I(\current_shift_inst.S3_syncZ0Z1 ));
    InMux I__6186 (
            .O(N__32246),
            .I(N__32240));
    InMux I__6185 (
            .O(N__32245),
            .I(N__32240));
    LocalMux I__6184 (
            .O(N__32240),
            .I(N__32236));
    InMux I__6183 (
            .O(N__32239),
            .I(N__32233));
    Span4Mux_h I__6182 (
            .O(N__32236),
            .I(N__32230));
    LocalMux I__6181 (
            .O(N__32233),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__6180 (
            .O(N__32230),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__6179 (
            .O(N__32225),
            .I(N__32222));
    LocalMux I__6178 (
            .O(N__32222),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ));
    InMux I__6177 (
            .O(N__32219),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__6176 (
            .O(N__32216),
            .I(N__32212));
    CascadeMux I__6175 (
            .O(N__32215),
            .I(N__32209));
    InMux I__6174 (
            .O(N__32212),
            .I(N__32204));
    InMux I__6173 (
            .O(N__32209),
            .I(N__32204));
    LocalMux I__6172 (
            .O(N__32204),
            .I(N__32200));
    InMux I__6171 (
            .O(N__32203),
            .I(N__32197));
    Span4Mux_h I__6170 (
            .O(N__32200),
            .I(N__32194));
    LocalMux I__6169 (
            .O(N__32197),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__6168 (
            .O(N__32194),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__6167 (
            .O(N__32189),
            .I(N__32186));
    LocalMux I__6166 (
            .O(N__32186),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ));
    InMux I__6165 (
            .O(N__32183),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__6164 (
            .O(N__32180),
            .I(N__32176));
    CascadeMux I__6163 (
            .O(N__32179),
            .I(N__32173));
    InMux I__6162 (
            .O(N__32176),
            .I(N__32168));
    InMux I__6161 (
            .O(N__32173),
            .I(N__32168));
    LocalMux I__6160 (
            .O(N__32168),
            .I(N__32164));
    InMux I__6159 (
            .O(N__32167),
            .I(N__32161));
    Span4Mux_h I__6158 (
            .O(N__32164),
            .I(N__32158));
    LocalMux I__6157 (
            .O(N__32161),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__6156 (
            .O(N__32158),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__6155 (
            .O(N__32153),
            .I(N__32150));
    LocalMux I__6154 (
            .O(N__32150),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ));
    InMux I__6153 (
            .O(N__32147),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__6152 (
            .O(N__32144),
            .I(N__32140));
    InMux I__6151 (
            .O(N__32143),
            .I(N__32137));
    LocalMux I__6150 (
            .O(N__32140),
            .I(N__32133));
    LocalMux I__6149 (
            .O(N__32137),
            .I(N__32130));
    InMux I__6148 (
            .O(N__32136),
            .I(N__32127));
    Span4Mux_h I__6147 (
            .O(N__32133),
            .I(N__32124));
    Span4Mux_h I__6146 (
            .O(N__32130),
            .I(N__32121));
    LocalMux I__6145 (
            .O(N__32127),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__6144 (
            .O(N__32124),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__6143 (
            .O(N__32121),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__6142 (
            .O(N__32114),
            .I(N__32111));
    LocalMux I__6141 (
            .O(N__32111),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ));
    InMux I__6140 (
            .O(N__32108),
            .I(bfn_12_22_0_));
    InMux I__6139 (
            .O(N__32105),
            .I(N__32101));
    InMux I__6138 (
            .O(N__32104),
            .I(N__32098));
    LocalMux I__6137 (
            .O(N__32101),
            .I(N__32094));
    LocalMux I__6136 (
            .O(N__32098),
            .I(N__32091));
    InMux I__6135 (
            .O(N__32097),
            .I(N__32088));
    Span4Mux_h I__6134 (
            .O(N__32094),
            .I(N__32085));
    Span4Mux_h I__6133 (
            .O(N__32091),
            .I(N__32082));
    LocalMux I__6132 (
            .O(N__32088),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__6131 (
            .O(N__32085),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__6130 (
            .O(N__32082),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__6129 (
            .O(N__32075),
            .I(N__32072));
    LocalMux I__6128 (
            .O(N__32072),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ));
    InMux I__6127 (
            .O(N__32069),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__6126 (
            .O(N__32066),
            .I(N__32063));
    LocalMux I__6125 (
            .O(N__32063),
            .I(N__32059));
    InMux I__6124 (
            .O(N__32062),
            .I(N__32056));
    Span4Mux_h I__6123 (
            .O(N__32059),
            .I(N__32053));
    LocalMux I__6122 (
            .O(N__32056),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__6121 (
            .O(N__32053),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    CascadeMux I__6120 (
            .O(N__32048),
            .I(N__32044));
    CascadeMux I__6119 (
            .O(N__32047),
            .I(N__32041));
    InMux I__6118 (
            .O(N__32044),
            .I(N__32035));
    InMux I__6117 (
            .O(N__32041),
            .I(N__32035));
    InMux I__6116 (
            .O(N__32040),
            .I(N__32032));
    LocalMux I__6115 (
            .O(N__32035),
            .I(N__32029));
    LocalMux I__6114 (
            .O(N__32032),
            .I(N__32024));
    Span4Mux_v I__6113 (
            .O(N__32029),
            .I(N__32024));
    Odrv4 I__6112 (
            .O(N__32024),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__6111 (
            .O(N__32021),
            .I(N__32018));
    LocalMux I__6110 (
            .O(N__32018),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ));
    InMux I__6109 (
            .O(N__32015),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__6108 (
            .O(N__32012),
            .I(N__32009));
    LocalMux I__6107 (
            .O(N__32009),
            .I(N__32005));
    InMux I__6106 (
            .O(N__32008),
            .I(N__32002));
    Span4Mux_h I__6105 (
            .O(N__32005),
            .I(N__31999));
    LocalMux I__6104 (
            .O(N__32002),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__6103 (
            .O(N__31999),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CascadeMux I__6102 (
            .O(N__31994),
            .I(N__31990));
    CascadeMux I__6101 (
            .O(N__31993),
            .I(N__31987));
    InMux I__6100 (
            .O(N__31990),
            .I(N__31981));
    InMux I__6099 (
            .O(N__31987),
            .I(N__31981));
    InMux I__6098 (
            .O(N__31986),
            .I(N__31978));
    LocalMux I__6097 (
            .O(N__31981),
            .I(N__31975));
    LocalMux I__6096 (
            .O(N__31978),
            .I(N__31970));
    Span4Mux_v I__6095 (
            .O(N__31975),
            .I(N__31970));
    Odrv4 I__6094 (
            .O(N__31970),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__6093 (
            .O(N__31967),
            .I(N__31964));
    LocalMux I__6092 (
            .O(N__31964),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ));
    InMux I__6091 (
            .O(N__31961),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__6090 (
            .O(N__31958),
            .I(N__31940));
    CEMux I__6089 (
            .O(N__31957),
            .I(N__31940));
    CEMux I__6088 (
            .O(N__31956),
            .I(N__31940));
    CEMux I__6087 (
            .O(N__31955),
            .I(N__31940));
    CEMux I__6086 (
            .O(N__31954),
            .I(N__31940));
    CEMux I__6085 (
            .O(N__31953),
            .I(N__31940));
    GlobalMux I__6084 (
            .O(N__31940),
            .I(N__31937));
    gio2CtrlBuf I__6083 (
            .O(N__31937),
            .I(\current_shift_inst.timer_s1.N_187_i_g ));
    InMux I__6082 (
            .O(N__31934),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__6081 (
            .O(N__31931),
            .I(N__31928));
    LocalMux I__6080 (
            .O(N__31928),
            .I(N__31924));
    InMux I__6079 (
            .O(N__31927),
            .I(N__31921));
    Span4Mux_h I__6078 (
            .O(N__31924),
            .I(N__31918));
    LocalMux I__6077 (
            .O(N__31921),
            .I(N__31915));
    Span4Mux_h I__6076 (
            .O(N__31918),
            .I(N__31910));
    Span4Mux_v I__6075 (
            .O(N__31915),
            .I(N__31910));
    Odrv4 I__6074 (
            .O(N__31910),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__6073 (
            .O(N__31907),
            .I(N__31901));
    InMux I__6072 (
            .O(N__31906),
            .I(N__31901));
    LocalMux I__6071 (
            .O(N__31901),
            .I(N__31897));
    InMux I__6070 (
            .O(N__31900),
            .I(N__31894));
    Span4Mux_h I__6069 (
            .O(N__31897),
            .I(N__31891));
    LocalMux I__6068 (
            .O(N__31894),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__6067 (
            .O(N__31891),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__6066 (
            .O(N__31886),
            .I(N__31883));
    LocalMux I__6065 (
            .O(N__31883),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ));
    InMux I__6064 (
            .O(N__31880),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__6063 (
            .O(N__31877),
            .I(N__31873));
    CascadeMux I__6062 (
            .O(N__31876),
            .I(N__31870));
    InMux I__6061 (
            .O(N__31873),
            .I(N__31865));
    InMux I__6060 (
            .O(N__31870),
            .I(N__31865));
    LocalMux I__6059 (
            .O(N__31865),
            .I(N__31861));
    InMux I__6058 (
            .O(N__31864),
            .I(N__31858));
    Span4Mux_h I__6057 (
            .O(N__31861),
            .I(N__31855));
    LocalMux I__6056 (
            .O(N__31858),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__6055 (
            .O(N__31855),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__6054 (
            .O(N__31850),
            .I(N__31847));
    LocalMux I__6053 (
            .O(N__31847),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ));
    InMux I__6052 (
            .O(N__31844),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__6051 (
            .O(N__31841),
            .I(N__31837));
    CascadeMux I__6050 (
            .O(N__31840),
            .I(N__31834));
    InMux I__6049 (
            .O(N__31837),
            .I(N__31829));
    InMux I__6048 (
            .O(N__31834),
            .I(N__31829));
    LocalMux I__6047 (
            .O(N__31829),
            .I(N__31825));
    InMux I__6046 (
            .O(N__31828),
            .I(N__31822));
    Span4Mux_h I__6045 (
            .O(N__31825),
            .I(N__31819));
    LocalMux I__6044 (
            .O(N__31822),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__6043 (
            .O(N__31819),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__6042 (
            .O(N__31814),
            .I(N__31811));
    LocalMux I__6041 (
            .O(N__31811),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ));
    InMux I__6040 (
            .O(N__31808),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__6039 (
            .O(N__31805),
            .I(N__31801));
    InMux I__6038 (
            .O(N__31804),
            .I(N__31798));
    LocalMux I__6037 (
            .O(N__31801),
            .I(N__31794));
    LocalMux I__6036 (
            .O(N__31798),
            .I(N__31791));
    InMux I__6035 (
            .O(N__31797),
            .I(N__31788));
    Span4Mux_h I__6034 (
            .O(N__31794),
            .I(N__31785));
    Span4Mux_h I__6033 (
            .O(N__31791),
            .I(N__31782));
    LocalMux I__6032 (
            .O(N__31788),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__6031 (
            .O(N__31785),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__6030 (
            .O(N__31782),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__6029 (
            .O(N__31775),
            .I(N__31772));
    LocalMux I__6028 (
            .O(N__31772),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ));
    InMux I__6027 (
            .O(N__31769),
            .I(bfn_12_21_0_));
    InMux I__6026 (
            .O(N__31766),
            .I(N__31762));
    InMux I__6025 (
            .O(N__31765),
            .I(N__31759));
    LocalMux I__6024 (
            .O(N__31762),
            .I(N__31755));
    LocalMux I__6023 (
            .O(N__31759),
            .I(N__31752));
    InMux I__6022 (
            .O(N__31758),
            .I(N__31749));
    Span4Mux_h I__6021 (
            .O(N__31755),
            .I(N__31746));
    Span4Mux_h I__6020 (
            .O(N__31752),
            .I(N__31743));
    LocalMux I__6019 (
            .O(N__31749),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__6018 (
            .O(N__31746),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__6017 (
            .O(N__31743),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__6016 (
            .O(N__31736),
            .I(N__31733));
    LocalMux I__6015 (
            .O(N__31733),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ));
    InMux I__6014 (
            .O(N__31730),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__6013 (
            .O(N__31727),
            .I(N__31723));
    CascadeMux I__6012 (
            .O(N__31726),
            .I(N__31720));
    InMux I__6011 (
            .O(N__31723),
            .I(N__31714));
    InMux I__6010 (
            .O(N__31720),
            .I(N__31714));
    InMux I__6009 (
            .O(N__31719),
            .I(N__31711));
    LocalMux I__6008 (
            .O(N__31714),
            .I(N__31708));
    LocalMux I__6007 (
            .O(N__31711),
            .I(N__31703));
    Span4Mux_v I__6006 (
            .O(N__31708),
            .I(N__31703));
    Odrv4 I__6005 (
            .O(N__31703),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__6004 (
            .O(N__31700),
            .I(N__31697));
    LocalMux I__6003 (
            .O(N__31697),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ));
    InMux I__6002 (
            .O(N__31694),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__6001 (
            .O(N__31691),
            .I(N__31687));
    CascadeMux I__6000 (
            .O(N__31690),
            .I(N__31684));
    InMux I__5999 (
            .O(N__31687),
            .I(N__31678));
    InMux I__5998 (
            .O(N__31684),
            .I(N__31678));
    InMux I__5997 (
            .O(N__31683),
            .I(N__31675));
    LocalMux I__5996 (
            .O(N__31678),
            .I(N__31672));
    LocalMux I__5995 (
            .O(N__31675),
            .I(N__31667));
    Span4Mux_v I__5994 (
            .O(N__31672),
            .I(N__31667));
    Odrv4 I__5993 (
            .O(N__31667),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__5992 (
            .O(N__31664),
            .I(N__31661));
    LocalMux I__5991 (
            .O(N__31661),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ));
    InMux I__5990 (
            .O(N__31658),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__5989 (
            .O(N__31655),
            .I(N__31649));
    InMux I__5988 (
            .O(N__31654),
            .I(N__31649));
    LocalMux I__5987 (
            .O(N__31649),
            .I(N__31645));
    InMux I__5986 (
            .O(N__31648),
            .I(N__31642));
    Span4Mux_h I__5985 (
            .O(N__31645),
            .I(N__31639));
    LocalMux I__5984 (
            .O(N__31642),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__5983 (
            .O(N__31639),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__5982 (
            .O(N__31634),
            .I(N__31631));
    LocalMux I__5981 (
            .O(N__31631),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ));
    InMux I__5980 (
            .O(N__31628),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__5979 (
            .O(N__31625),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__5978 (
            .O(N__31622),
            .I(N__31616));
    InMux I__5977 (
            .O(N__31621),
            .I(N__31616));
    LocalMux I__5976 (
            .O(N__31616),
            .I(N__31612));
    InMux I__5975 (
            .O(N__31615),
            .I(N__31609));
    Span4Mux_h I__5974 (
            .O(N__31612),
            .I(N__31606));
    LocalMux I__5973 (
            .O(N__31609),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__5972 (
            .O(N__31606),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__5971 (
            .O(N__31601),
            .I(N__31598));
    LocalMux I__5970 (
            .O(N__31598),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ));
    InMux I__5969 (
            .O(N__31595),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__5968 (
            .O(N__31592),
            .I(N__31586));
    InMux I__5967 (
            .O(N__31591),
            .I(N__31586));
    LocalMux I__5966 (
            .O(N__31586),
            .I(N__31582));
    InMux I__5965 (
            .O(N__31585),
            .I(N__31579));
    Span4Mux_h I__5964 (
            .O(N__31582),
            .I(N__31576));
    LocalMux I__5963 (
            .O(N__31579),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__5962 (
            .O(N__31576),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__5961 (
            .O(N__31571),
            .I(N__31568));
    LocalMux I__5960 (
            .O(N__31568),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ));
    InMux I__5959 (
            .O(N__31565),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__5958 (
            .O(N__31562),
            .I(N__31558));
    InMux I__5957 (
            .O(N__31561),
            .I(N__31555));
    InMux I__5956 (
            .O(N__31558),
            .I(N__31552));
    LocalMux I__5955 (
            .O(N__31555),
            .I(N__31548));
    LocalMux I__5954 (
            .O(N__31552),
            .I(N__31545));
    InMux I__5953 (
            .O(N__31551),
            .I(N__31542));
    Span4Mux_h I__5952 (
            .O(N__31548),
            .I(N__31539));
    Span4Mux_h I__5951 (
            .O(N__31545),
            .I(N__31536));
    LocalMux I__5950 (
            .O(N__31542),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__5949 (
            .O(N__31539),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__5948 (
            .O(N__31536),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__5947 (
            .O(N__31529),
            .I(N__31526));
    LocalMux I__5946 (
            .O(N__31526),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ));
    InMux I__5945 (
            .O(N__31523),
            .I(bfn_12_20_0_));
    CascadeMux I__5944 (
            .O(N__31520),
            .I(N__31516));
    InMux I__5943 (
            .O(N__31519),
            .I(N__31513));
    InMux I__5942 (
            .O(N__31516),
            .I(N__31510));
    LocalMux I__5941 (
            .O(N__31513),
            .I(N__31506));
    LocalMux I__5940 (
            .O(N__31510),
            .I(N__31503));
    InMux I__5939 (
            .O(N__31509),
            .I(N__31500));
    Span4Mux_h I__5938 (
            .O(N__31506),
            .I(N__31497));
    Span4Mux_h I__5937 (
            .O(N__31503),
            .I(N__31494));
    LocalMux I__5936 (
            .O(N__31500),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__5935 (
            .O(N__31497),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__5934 (
            .O(N__31494),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__5933 (
            .O(N__31487),
            .I(N__31484));
    LocalMux I__5932 (
            .O(N__31484),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ));
    InMux I__5931 (
            .O(N__31481),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__5930 (
            .O(N__31478),
            .I(N__31474));
    CascadeMux I__5929 (
            .O(N__31477),
            .I(N__31471));
    InMux I__5928 (
            .O(N__31474),
            .I(N__31465));
    InMux I__5927 (
            .O(N__31471),
            .I(N__31465));
    InMux I__5926 (
            .O(N__31470),
            .I(N__31462));
    LocalMux I__5925 (
            .O(N__31465),
            .I(N__31459));
    LocalMux I__5924 (
            .O(N__31462),
            .I(N__31454));
    Span4Mux_v I__5923 (
            .O(N__31459),
            .I(N__31454));
    Odrv4 I__5922 (
            .O(N__31454),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__5921 (
            .O(N__31451),
            .I(N__31448));
    LocalMux I__5920 (
            .O(N__31448),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ));
    InMux I__5919 (
            .O(N__31445),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__5918 (
            .O(N__31442),
            .I(N__31438));
    CascadeMux I__5917 (
            .O(N__31441),
            .I(N__31435));
    InMux I__5916 (
            .O(N__31438),
            .I(N__31429));
    InMux I__5915 (
            .O(N__31435),
            .I(N__31429));
    InMux I__5914 (
            .O(N__31434),
            .I(N__31426));
    LocalMux I__5913 (
            .O(N__31429),
            .I(N__31423));
    LocalMux I__5912 (
            .O(N__31426),
            .I(N__31418));
    Span4Mux_v I__5911 (
            .O(N__31423),
            .I(N__31418));
    Odrv4 I__5910 (
            .O(N__31418),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__5909 (
            .O(N__31415),
            .I(N__31412));
    LocalMux I__5908 (
            .O(N__31412),
            .I(N__31409));
    Odrv4 I__5907 (
            .O(N__31409),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ));
    InMux I__5906 (
            .O(N__31406),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__5905 (
            .O(N__31403),
            .I(N__31397));
    InMux I__5904 (
            .O(N__31402),
            .I(N__31397));
    LocalMux I__5903 (
            .O(N__31397),
            .I(N__31393));
    InMux I__5902 (
            .O(N__31396),
            .I(N__31390));
    Span4Mux_h I__5901 (
            .O(N__31393),
            .I(N__31387));
    LocalMux I__5900 (
            .O(N__31390),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__5899 (
            .O(N__31387),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__5898 (
            .O(N__31382),
            .I(N__31379));
    LocalMux I__5897 (
            .O(N__31379),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ));
    InMux I__5896 (
            .O(N__31376),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__5895 (
            .O(N__31373),
            .I(N__31367));
    InMux I__5894 (
            .O(N__31372),
            .I(N__31367));
    LocalMux I__5893 (
            .O(N__31367),
            .I(N__31363));
    InMux I__5892 (
            .O(N__31366),
            .I(N__31360));
    Span4Mux_h I__5891 (
            .O(N__31363),
            .I(N__31357));
    LocalMux I__5890 (
            .O(N__31360),
            .I(N__31354));
    Span4Mux_v I__5889 (
            .O(N__31357),
            .I(N__31350));
    Span4Mux_v I__5888 (
            .O(N__31354),
            .I(N__31347));
    InMux I__5887 (
            .O(N__31353),
            .I(N__31344));
    Odrv4 I__5886 (
            .O(N__31350),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    Odrv4 I__5885 (
            .O(N__31347),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    LocalMux I__5884 (
            .O(N__31344),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    CascadeMux I__5883 (
            .O(N__31337),
            .I(N__31333));
    InMux I__5882 (
            .O(N__31336),
            .I(N__31329));
    InMux I__5881 (
            .O(N__31333),
            .I(N__31324));
    InMux I__5880 (
            .O(N__31332),
            .I(N__31324));
    LocalMux I__5879 (
            .O(N__31329),
            .I(N__31320));
    LocalMux I__5878 (
            .O(N__31324),
            .I(N__31317));
    CascadeMux I__5877 (
            .O(N__31323),
            .I(N__31314));
    Span4Mux_h I__5876 (
            .O(N__31320),
            .I(N__31311));
    Span4Mux_h I__5875 (
            .O(N__31317),
            .I(N__31308));
    InMux I__5874 (
            .O(N__31314),
            .I(N__31305));
    Odrv4 I__5873 (
            .O(N__31311),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    Odrv4 I__5872 (
            .O(N__31308),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    LocalMux I__5871 (
            .O(N__31305),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    CascadeMux I__5870 (
            .O(N__31298),
            .I(N__31295));
    InMux I__5869 (
            .O(N__31295),
            .I(N__31292));
    LocalMux I__5868 (
            .O(N__31292),
            .I(N__31289));
    Span4Mux_h I__5867 (
            .O(N__31289),
            .I(N__31286));
    Odrv4 I__5866 (
            .O(N__31286),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ));
    InMux I__5865 (
            .O(N__31283),
            .I(N__31279));
    InMux I__5864 (
            .O(N__31282),
            .I(N__31276));
    LocalMux I__5863 (
            .O(N__31279),
            .I(N__31272));
    LocalMux I__5862 (
            .O(N__31276),
            .I(N__31268));
    CascadeMux I__5861 (
            .O(N__31275),
            .I(N__31265));
    Span4Mux_h I__5860 (
            .O(N__31272),
            .I(N__31262));
    InMux I__5859 (
            .O(N__31271),
            .I(N__31259));
    Span4Mux_v I__5858 (
            .O(N__31268),
            .I(N__31256));
    InMux I__5857 (
            .O(N__31265),
            .I(N__31253));
    Span4Mux_h I__5856 (
            .O(N__31262),
            .I(N__31250));
    LocalMux I__5855 (
            .O(N__31259),
            .I(N__31247));
    Span4Mux_h I__5854 (
            .O(N__31256),
            .I(N__31242));
    LocalMux I__5853 (
            .O(N__31253),
            .I(N__31242));
    Odrv4 I__5852 (
            .O(N__31250),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    Odrv12 I__5851 (
            .O(N__31247),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    Odrv4 I__5850 (
            .O(N__31242),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    CascadeMux I__5849 (
            .O(N__31235),
            .I(N__31232));
    InMux I__5848 (
            .O(N__31232),
            .I(N__31227));
    InMux I__5847 (
            .O(N__31231),
            .I(N__31224));
    InMux I__5846 (
            .O(N__31230),
            .I(N__31221));
    LocalMux I__5845 (
            .O(N__31227),
            .I(N__31215));
    LocalMux I__5844 (
            .O(N__31224),
            .I(N__31215));
    LocalMux I__5843 (
            .O(N__31221),
            .I(N__31212));
    CascadeMux I__5842 (
            .O(N__31220),
            .I(N__31209));
    Span4Mux_h I__5841 (
            .O(N__31215),
            .I(N__31206));
    Span4Mux_h I__5840 (
            .O(N__31212),
            .I(N__31203));
    InMux I__5839 (
            .O(N__31209),
            .I(N__31200));
    Odrv4 I__5838 (
            .O(N__31206),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    Odrv4 I__5837 (
            .O(N__31203),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    LocalMux I__5836 (
            .O(N__31200),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    CascadeMux I__5835 (
            .O(N__31193),
            .I(N__31190));
    InMux I__5834 (
            .O(N__31190),
            .I(N__31185));
    InMux I__5833 (
            .O(N__31189),
            .I(N__31182));
    InMux I__5832 (
            .O(N__31188),
            .I(N__31179));
    LocalMux I__5831 (
            .O(N__31185),
            .I(N__31175));
    LocalMux I__5830 (
            .O(N__31182),
            .I(N__31172));
    LocalMux I__5829 (
            .O(N__31179),
            .I(N__31169));
    CascadeMux I__5828 (
            .O(N__31178),
            .I(N__31166));
    Span4Mux_v I__5827 (
            .O(N__31175),
            .I(N__31163));
    Span4Mux_h I__5826 (
            .O(N__31172),
            .I(N__31160));
    Span4Mux_h I__5825 (
            .O(N__31169),
            .I(N__31157));
    InMux I__5824 (
            .O(N__31166),
            .I(N__31154));
    Odrv4 I__5823 (
            .O(N__31163),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    Odrv4 I__5822 (
            .O(N__31160),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    Odrv4 I__5821 (
            .O(N__31157),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    LocalMux I__5820 (
            .O(N__31154),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    InMux I__5819 (
            .O(N__31145),
            .I(N__31142));
    LocalMux I__5818 (
            .O(N__31142),
            .I(N__31137));
    InMux I__5817 (
            .O(N__31141),
            .I(N__31132));
    InMux I__5816 (
            .O(N__31140),
            .I(N__31132));
    Span4Mux_h I__5815 (
            .O(N__31137),
            .I(N__31129));
    LocalMux I__5814 (
            .O(N__31132),
            .I(N__31125));
    Span4Mux_h I__5813 (
            .O(N__31129),
            .I(N__31122));
    InMux I__5812 (
            .O(N__31128),
            .I(N__31119));
    Odrv12 I__5811 (
            .O(N__31125),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    Odrv4 I__5810 (
            .O(N__31122),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    LocalMux I__5809 (
            .O(N__31119),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    InMux I__5808 (
            .O(N__31112),
            .I(N__31109));
    LocalMux I__5807 (
            .O(N__31109),
            .I(N__31106));
    Span4Mux_h I__5806 (
            .O(N__31106),
            .I(N__31103));
    Odrv4 I__5805 (
            .O(N__31103),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ));
    CascadeMux I__5804 (
            .O(N__31100),
            .I(N__31096));
    InMux I__5803 (
            .O(N__31099),
            .I(N__31093));
    InMux I__5802 (
            .O(N__31096),
            .I(N__31090));
    LocalMux I__5801 (
            .O(N__31093),
            .I(N__31087));
    LocalMux I__5800 (
            .O(N__31090),
            .I(N__31083));
    Span4Mux_v I__5799 (
            .O(N__31087),
            .I(N__31080));
    InMux I__5798 (
            .O(N__31086),
            .I(N__31077));
    Span4Mux_h I__5797 (
            .O(N__31083),
            .I(N__31074));
    Odrv4 I__5796 (
            .O(N__31080),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__5795 (
            .O(N__31077),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__5794 (
            .O(N__31074),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__5793 (
            .O(N__31067),
            .I(N__31064));
    LocalMux I__5792 (
            .O(N__31064),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ));
    CascadeMux I__5791 (
            .O(N__31061),
            .I(N__31057));
    InMux I__5790 (
            .O(N__31060),
            .I(N__31054));
    InMux I__5789 (
            .O(N__31057),
            .I(N__31051));
    LocalMux I__5788 (
            .O(N__31054),
            .I(N__31048));
    LocalMux I__5787 (
            .O(N__31051),
            .I(N__31044));
    Span4Mux_v I__5786 (
            .O(N__31048),
            .I(N__31041));
    InMux I__5785 (
            .O(N__31047),
            .I(N__31038));
    Span4Mux_h I__5784 (
            .O(N__31044),
            .I(N__31035));
    Odrv4 I__5783 (
            .O(N__31041),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__5782 (
            .O(N__31038),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__5781 (
            .O(N__31035),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__5780 (
            .O(N__31028),
            .I(N__31025));
    LocalMux I__5779 (
            .O(N__31025),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ));
    InMux I__5778 (
            .O(N__31022),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__5777 (
            .O(N__31019),
            .I(N__31012));
    InMux I__5776 (
            .O(N__31018),
            .I(N__31012));
    InMux I__5775 (
            .O(N__31017),
            .I(N__31009));
    LocalMux I__5774 (
            .O(N__31012),
            .I(N__31006));
    LocalMux I__5773 (
            .O(N__31009),
            .I(N__31001));
    Span4Mux_v I__5772 (
            .O(N__31006),
            .I(N__31001));
    Odrv4 I__5771 (
            .O(N__31001),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__5770 (
            .O(N__30998),
            .I(N__30995));
    LocalMux I__5769 (
            .O(N__30995),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ));
    InMux I__5768 (
            .O(N__30992),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__5767 (
            .O(N__30989),
            .I(N__30982));
    InMux I__5766 (
            .O(N__30988),
            .I(N__30982));
    InMux I__5765 (
            .O(N__30987),
            .I(N__30979));
    LocalMux I__5764 (
            .O(N__30982),
            .I(N__30976));
    LocalMux I__5763 (
            .O(N__30979),
            .I(N__30971));
    Span4Mux_v I__5762 (
            .O(N__30976),
            .I(N__30971));
    Odrv4 I__5761 (
            .O(N__30971),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__5760 (
            .O(N__30968),
            .I(N__30965));
    LocalMux I__5759 (
            .O(N__30965),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ));
    InMux I__5758 (
            .O(N__30962),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__5757 (
            .O(N__30959),
            .I(N__30955));
    CascadeMux I__5756 (
            .O(N__30958),
            .I(N__30952));
    InMux I__5755 (
            .O(N__30955),
            .I(N__30947));
    InMux I__5754 (
            .O(N__30952),
            .I(N__30947));
    LocalMux I__5753 (
            .O(N__30947),
            .I(N__30943));
    InMux I__5752 (
            .O(N__30946),
            .I(N__30940));
    Span4Mux_h I__5751 (
            .O(N__30943),
            .I(N__30937));
    LocalMux I__5750 (
            .O(N__30940),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__5749 (
            .O(N__30937),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__5748 (
            .O(N__30932),
            .I(N__30929));
    LocalMux I__5747 (
            .O(N__30929),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ));
    InMux I__5746 (
            .O(N__30926),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__5745 (
            .O(N__30923),
            .I(N__30919));
    CascadeMux I__5744 (
            .O(N__30922),
            .I(N__30916));
    InMux I__5743 (
            .O(N__30919),
            .I(N__30911));
    InMux I__5742 (
            .O(N__30916),
            .I(N__30911));
    LocalMux I__5741 (
            .O(N__30911),
            .I(N__30907));
    InMux I__5740 (
            .O(N__30910),
            .I(N__30904));
    Span4Mux_h I__5739 (
            .O(N__30907),
            .I(N__30901));
    LocalMux I__5738 (
            .O(N__30904),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__5737 (
            .O(N__30901),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__5736 (
            .O(N__30896),
            .I(N__30893));
    LocalMux I__5735 (
            .O(N__30893),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ));
    InMux I__5734 (
            .O(N__30890),
            .I(N__30887));
    LocalMux I__5733 (
            .O(N__30887),
            .I(N__30882));
    InMux I__5732 (
            .O(N__30886),
            .I(N__30879));
    InMux I__5731 (
            .O(N__30885),
            .I(N__30876));
    Span4Mux_v I__5730 (
            .O(N__30882),
            .I(N__30871));
    LocalMux I__5729 (
            .O(N__30879),
            .I(N__30871));
    LocalMux I__5728 (
            .O(N__30876),
            .I(N__30868));
    Span4Mux_h I__5727 (
            .O(N__30871),
            .I(N__30864));
    Span4Mux_h I__5726 (
            .O(N__30868),
            .I(N__30861));
    InMux I__5725 (
            .O(N__30867),
            .I(N__30858));
    Span4Mux_v I__5724 (
            .O(N__30864),
            .I(N__30855));
    Span4Mux_h I__5723 (
            .O(N__30861),
            .I(N__30850));
    LocalMux I__5722 (
            .O(N__30858),
            .I(N__30850));
    Odrv4 I__5721 (
            .O(N__30855),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    Odrv4 I__5720 (
            .O(N__30850),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    InMux I__5719 (
            .O(N__30845),
            .I(N__30840));
    InMux I__5718 (
            .O(N__30844),
            .I(N__30837));
    InMux I__5717 (
            .O(N__30843),
            .I(N__30834));
    LocalMux I__5716 (
            .O(N__30840),
            .I(N__30831));
    LocalMux I__5715 (
            .O(N__30837),
            .I(N__30828));
    LocalMux I__5714 (
            .O(N__30834),
            .I(N__30824));
    Span4Mux_h I__5713 (
            .O(N__30831),
            .I(N__30819));
    Span4Mux_h I__5712 (
            .O(N__30828),
            .I(N__30819));
    InMux I__5711 (
            .O(N__30827),
            .I(N__30816));
    Odrv12 I__5710 (
            .O(N__30824),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    Odrv4 I__5709 (
            .O(N__30819),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    LocalMux I__5708 (
            .O(N__30816),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    CascadeMux I__5707 (
            .O(N__30809),
            .I(N__30806));
    InMux I__5706 (
            .O(N__30806),
            .I(N__30802));
    InMux I__5705 (
            .O(N__30805),
            .I(N__30798));
    LocalMux I__5704 (
            .O(N__30802),
            .I(N__30794));
    InMux I__5703 (
            .O(N__30801),
            .I(N__30791));
    LocalMux I__5702 (
            .O(N__30798),
            .I(N__30788));
    CascadeMux I__5701 (
            .O(N__30797),
            .I(N__30785));
    Span4Mux_h I__5700 (
            .O(N__30794),
            .I(N__30782));
    LocalMux I__5699 (
            .O(N__30791),
            .I(N__30779));
    Span4Mux_h I__5698 (
            .O(N__30788),
            .I(N__30776));
    InMux I__5697 (
            .O(N__30785),
            .I(N__30773));
    Odrv4 I__5696 (
            .O(N__30782),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    Odrv12 I__5695 (
            .O(N__30779),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    Odrv4 I__5694 (
            .O(N__30776),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    LocalMux I__5693 (
            .O(N__30773),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    InMux I__5692 (
            .O(N__30764),
            .I(N__30759));
    InMux I__5691 (
            .O(N__30763),
            .I(N__30756));
    InMux I__5690 (
            .O(N__30762),
            .I(N__30753));
    LocalMux I__5689 (
            .O(N__30759),
            .I(N__30750));
    LocalMux I__5688 (
            .O(N__30756),
            .I(N__30747));
    LocalMux I__5687 (
            .O(N__30753),
            .I(N__30741));
    Span4Mux_h I__5686 (
            .O(N__30750),
            .I(N__30741));
    Span4Mux_h I__5685 (
            .O(N__30747),
            .I(N__30738));
    InMux I__5684 (
            .O(N__30746),
            .I(N__30735));
    Span4Mux_v I__5683 (
            .O(N__30741),
            .I(N__30728));
    Span4Mux_h I__5682 (
            .O(N__30738),
            .I(N__30728));
    LocalMux I__5681 (
            .O(N__30735),
            .I(N__30728));
    Odrv4 I__5680 (
            .O(N__30728),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    InMux I__5679 (
            .O(N__30725),
            .I(N__30722));
    LocalMux I__5678 (
            .O(N__30722),
            .I(N__30719));
    Span4Mux_h I__5677 (
            .O(N__30719),
            .I(N__30716));
    Odrv4 I__5676 (
            .O(N__30716),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ));
    CascadeMux I__5675 (
            .O(N__30713),
            .I(N__30710));
    InMux I__5674 (
            .O(N__30710),
            .I(N__30707));
    LocalMux I__5673 (
            .O(N__30707),
            .I(N__30704));
    Span4Mux_h I__5672 (
            .O(N__30704),
            .I(N__30701));
    Odrv4 I__5671 (
            .O(N__30701),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ));
    InMux I__5670 (
            .O(N__30698),
            .I(N__30693));
    InMux I__5669 (
            .O(N__30697),
            .I(N__30690));
    InMux I__5668 (
            .O(N__30696),
            .I(N__30687));
    LocalMux I__5667 (
            .O(N__30693),
            .I(N__30684));
    LocalMux I__5666 (
            .O(N__30690),
            .I(N__30680));
    LocalMux I__5665 (
            .O(N__30687),
            .I(N__30677));
    Span4Mux_v I__5664 (
            .O(N__30684),
            .I(N__30674));
    InMux I__5663 (
            .O(N__30683),
            .I(N__30671));
    Span4Mux_v I__5662 (
            .O(N__30680),
            .I(N__30668));
    Span4Mux_v I__5661 (
            .O(N__30677),
            .I(N__30661));
    Span4Mux_h I__5660 (
            .O(N__30674),
            .I(N__30661));
    LocalMux I__5659 (
            .O(N__30671),
            .I(N__30661));
    Odrv4 I__5658 (
            .O(N__30668),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    Odrv4 I__5657 (
            .O(N__30661),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    InMux I__5656 (
            .O(N__30656),
            .I(N__30651));
    CascadeMux I__5655 (
            .O(N__30655),
            .I(N__30648));
    InMux I__5654 (
            .O(N__30654),
            .I(N__30645));
    LocalMux I__5653 (
            .O(N__30651),
            .I(N__30641));
    InMux I__5652 (
            .O(N__30648),
            .I(N__30638));
    LocalMux I__5651 (
            .O(N__30645),
            .I(N__30635));
    CascadeMux I__5650 (
            .O(N__30644),
            .I(N__30632));
    Span4Mux_h I__5649 (
            .O(N__30641),
            .I(N__30629));
    LocalMux I__5648 (
            .O(N__30638),
            .I(N__30624));
    Span4Mux_h I__5647 (
            .O(N__30635),
            .I(N__30624));
    InMux I__5646 (
            .O(N__30632),
            .I(N__30621));
    Odrv4 I__5645 (
            .O(N__30629),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    Odrv4 I__5644 (
            .O(N__30624),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    LocalMux I__5643 (
            .O(N__30621),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    InMux I__5642 (
            .O(N__30614),
            .I(N__30611));
    LocalMux I__5641 (
            .O(N__30611),
            .I(N__30608));
    Span4Mux_h I__5640 (
            .O(N__30608),
            .I(N__30605));
    Odrv4 I__5639 (
            .O(N__30605),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ));
    InMux I__5638 (
            .O(N__30602),
            .I(N__30599));
    LocalMux I__5637 (
            .O(N__30599),
            .I(N__30593));
    CascadeMux I__5636 (
            .O(N__30598),
            .I(N__30590));
    InMux I__5635 (
            .O(N__30597),
            .I(N__30585));
    InMux I__5634 (
            .O(N__30596),
            .I(N__30585));
    Span4Mux_h I__5633 (
            .O(N__30593),
            .I(N__30582));
    InMux I__5632 (
            .O(N__30590),
            .I(N__30579));
    LocalMux I__5631 (
            .O(N__30585),
            .I(N__30576));
    Span4Mux_h I__5630 (
            .O(N__30582),
            .I(N__30571));
    LocalMux I__5629 (
            .O(N__30579),
            .I(N__30571));
    Odrv12 I__5628 (
            .O(N__30576),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    Odrv4 I__5627 (
            .O(N__30571),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    CascadeMux I__5626 (
            .O(N__30566),
            .I(N__30563));
    InMux I__5625 (
            .O(N__30563),
            .I(N__30556));
    InMux I__5624 (
            .O(N__30562),
            .I(N__30556));
    InMux I__5623 (
            .O(N__30561),
            .I(N__30553));
    LocalMux I__5622 (
            .O(N__30556),
            .I(N__30549));
    LocalMux I__5621 (
            .O(N__30553),
            .I(N__30546));
    CascadeMux I__5620 (
            .O(N__30552),
            .I(N__30543));
    Span4Mux_h I__5619 (
            .O(N__30549),
            .I(N__30540));
    Span4Mux_h I__5618 (
            .O(N__30546),
            .I(N__30537));
    InMux I__5617 (
            .O(N__30543),
            .I(N__30534));
    Odrv4 I__5616 (
            .O(N__30540),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    Odrv4 I__5615 (
            .O(N__30537),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    LocalMux I__5614 (
            .O(N__30534),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    InMux I__5613 (
            .O(N__30527),
            .I(N__30524));
    LocalMux I__5612 (
            .O(N__30524),
            .I(N__30521));
    Span4Mux_h I__5611 (
            .O(N__30521),
            .I(N__30518));
    Odrv4 I__5610 (
            .O(N__30518),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ));
    CascadeMux I__5609 (
            .O(N__30515),
            .I(N__30512));
    InMux I__5608 (
            .O(N__30512),
            .I(N__30509));
    LocalMux I__5607 (
            .O(N__30509),
            .I(N__30503));
    InMux I__5606 (
            .O(N__30508),
            .I(N__30498));
    InMux I__5605 (
            .O(N__30507),
            .I(N__30498));
    CascadeMux I__5604 (
            .O(N__30506),
            .I(N__30495));
    Span4Mux_v I__5603 (
            .O(N__30503),
            .I(N__30492));
    LocalMux I__5602 (
            .O(N__30498),
            .I(N__30489));
    InMux I__5601 (
            .O(N__30495),
            .I(N__30486));
    Span4Mux_h I__5600 (
            .O(N__30492),
            .I(N__30483));
    Span12Mux_v I__5599 (
            .O(N__30489),
            .I(N__30480));
    LocalMux I__5598 (
            .O(N__30486),
            .I(N__30477));
    Odrv4 I__5597 (
            .O(N__30483),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    Odrv12 I__5596 (
            .O(N__30480),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    Odrv4 I__5595 (
            .O(N__30477),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    CascadeMux I__5594 (
            .O(N__30470),
            .I(N__30467));
    InMux I__5593 (
            .O(N__30467),
            .I(N__30460));
    InMux I__5592 (
            .O(N__30466),
            .I(N__30460));
    InMux I__5591 (
            .O(N__30465),
            .I(N__30456));
    LocalMux I__5590 (
            .O(N__30460),
            .I(N__30453));
    CascadeMux I__5589 (
            .O(N__30459),
            .I(N__30450));
    LocalMux I__5588 (
            .O(N__30456),
            .I(N__30447));
    Span4Mux_h I__5587 (
            .O(N__30453),
            .I(N__30444));
    InMux I__5586 (
            .O(N__30450),
            .I(N__30441));
    Odrv12 I__5585 (
            .O(N__30447),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    Odrv4 I__5584 (
            .O(N__30444),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    LocalMux I__5583 (
            .O(N__30441),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    CascadeMux I__5582 (
            .O(N__30434),
            .I(N__30431));
    InMux I__5581 (
            .O(N__30431),
            .I(N__30428));
    LocalMux I__5580 (
            .O(N__30428),
            .I(N__30425));
    Span4Mux_v I__5579 (
            .O(N__30425),
            .I(N__30422));
    Odrv4 I__5578 (
            .O(N__30422),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ));
    CascadeMux I__5577 (
            .O(N__30419),
            .I(N__30416));
    InMux I__5576 (
            .O(N__30416),
            .I(N__30413));
    LocalMux I__5575 (
            .O(N__30413),
            .I(N__30410));
    Odrv4 I__5574 (
            .O(N__30410),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__5573 (
            .O(N__30407),
            .I(N__30404));
    InMux I__5572 (
            .O(N__30404),
            .I(N__30399));
    InMux I__5571 (
            .O(N__30403),
            .I(N__30396));
    CascadeMux I__5570 (
            .O(N__30402),
            .I(N__30393));
    LocalMux I__5569 (
            .O(N__30399),
            .I(N__30389));
    LocalMux I__5568 (
            .O(N__30396),
            .I(N__30386));
    InMux I__5567 (
            .O(N__30393),
            .I(N__30381));
    InMux I__5566 (
            .O(N__30392),
            .I(N__30381));
    Span12Mux_h I__5565 (
            .O(N__30389),
            .I(N__30378));
    Span4Mux_h I__5564 (
            .O(N__30386),
            .I(N__30375));
    LocalMux I__5563 (
            .O(N__30381),
            .I(N__30372));
    Odrv12 I__5562 (
            .O(N__30378),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__5561 (
            .O(N__30375),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__5560 (
            .O(N__30372),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__5559 (
            .O(N__30365),
            .I(N__30362));
    LocalMux I__5558 (
            .O(N__30362),
            .I(N__30359));
    Odrv4 I__5557 (
            .O(N__30359),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__5556 (
            .O(N__30356),
            .I(N__30353));
    LocalMux I__5555 (
            .O(N__30353),
            .I(N__30350));
    Span4Mux_h I__5554 (
            .O(N__30350),
            .I(N__30344));
    InMux I__5553 (
            .O(N__30349),
            .I(N__30341));
    InMux I__5552 (
            .O(N__30348),
            .I(N__30336));
    InMux I__5551 (
            .O(N__30347),
            .I(N__30336));
    Span4Mux_h I__5550 (
            .O(N__30344),
            .I(N__30333));
    LocalMux I__5549 (
            .O(N__30341),
            .I(N__30330));
    LocalMux I__5548 (
            .O(N__30336),
            .I(N__30327));
    Odrv4 I__5547 (
            .O(N__30333),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__5546 (
            .O(N__30330),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__5545 (
            .O(N__30327),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    CascadeMux I__5544 (
            .O(N__30320),
            .I(\phase_controller_inst1.stoper_hc.un1_m5_iZ0Z_1_cascade_ ));
    CascadeMux I__5543 (
            .O(N__30317),
            .I(\phase_controller_inst1.stoper_hc.un1_N_4_cascade_ ));
    InMux I__5542 (
            .O(N__30314),
            .I(N__30311));
    LocalMux I__5541 (
            .O(N__30311),
            .I(\current_shift_inst.S1_sync_prevZ0 ));
    InMux I__5540 (
            .O(N__30308),
            .I(N__30305));
    LocalMux I__5539 (
            .O(N__30305),
            .I(\current_shift_inst.S1_syncZ0Z0 ));
    InMux I__5538 (
            .O(N__30302),
            .I(N__30296));
    InMux I__5537 (
            .O(N__30301),
            .I(N__30296));
    LocalMux I__5536 (
            .O(N__30296),
            .I(\current_shift_inst.S1_syncZ0Z1 ));
    InMux I__5535 (
            .O(N__30293),
            .I(N__30290));
    LocalMux I__5534 (
            .O(N__30290),
            .I(N__30286));
    CascadeMux I__5533 (
            .O(N__30289),
            .I(N__30282));
    Span4Mux_h I__5532 (
            .O(N__30286),
            .I(N__30275));
    InMux I__5531 (
            .O(N__30285),
            .I(N__30272));
    InMux I__5530 (
            .O(N__30282),
            .I(N__30265));
    InMux I__5529 (
            .O(N__30281),
            .I(N__30265));
    InMux I__5528 (
            .O(N__30280),
            .I(N__30265));
    InMux I__5527 (
            .O(N__30279),
            .I(N__30262));
    InMux I__5526 (
            .O(N__30278),
            .I(N__30259));
    Odrv4 I__5525 (
            .O(N__30275),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__5524 (
            .O(N__30272),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__5523 (
            .O(N__30265),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__5522 (
            .O(N__30262),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__5521 (
            .O(N__30259),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    InMux I__5520 (
            .O(N__30248),
            .I(N__30237));
    InMux I__5519 (
            .O(N__30247),
            .I(N__30237));
    InMux I__5518 (
            .O(N__30246),
            .I(N__30237));
    InMux I__5517 (
            .O(N__30245),
            .I(N__30234));
    InMux I__5516 (
            .O(N__30244),
            .I(N__30229));
    LocalMux I__5515 (
            .O(N__30237),
            .I(N__30226));
    LocalMux I__5514 (
            .O(N__30234),
            .I(N__30223));
    InMux I__5513 (
            .O(N__30233),
            .I(N__30220));
    InMux I__5512 (
            .O(N__30232),
            .I(N__30217));
    LocalMux I__5511 (
            .O(N__30229),
            .I(N__30210));
    Span4Mux_v I__5510 (
            .O(N__30226),
            .I(N__30210));
    Span4Mux_v I__5509 (
            .O(N__30223),
            .I(N__30210));
    LocalMux I__5508 (
            .O(N__30220),
            .I(\current_shift_inst.S1_riseZ0 ));
    LocalMux I__5507 (
            .O(N__30217),
            .I(\current_shift_inst.S1_riseZ0 ));
    Odrv4 I__5506 (
            .O(N__30210),
            .I(\current_shift_inst.S1_riseZ0 ));
    InMux I__5505 (
            .O(N__30203),
            .I(N__30199));
    InMux I__5504 (
            .O(N__30202),
            .I(N__30195));
    LocalMux I__5503 (
            .O(N__30199),
            .I(N__30191));
    InMux I__5502 (
            .O(N__30198),
            .I(N__30188));
    LocalMux I__5501 (
            .O(N__30195),
            .I(N__30185));
    InMux I__5500 (
            .O(N__30194),
            .I(N__30181));
    Span12Mux_s8_h I__5499 (
            .O(N__30191),
            .I(N__30178));
    LocalMux I__5498 (
            .O(N__30188),
            .I(N__30175));
    Span4Mux_h I__5497 (
            .O(N__30185),
            .I(N__30172));
    InMux I__5496 (
            .O(N__30184),
            .I(N__30169));
    LocalMux I__5495 (
            .O(N__30181),
            .I(N__30164));
    Span12Mux_v I__5494 (
            .O(N__30178),
            .I(N__30164));
    Span4Mux_h I__5493 (
            .O(N__30175),
            .I(N__30161));
    Odrv4 I__5492 (
            .O(N__30172),
            .I(\current_shift_inst.phase_validZ0 ));
    LocalMux I__5491 (
            .O(N__30169),
            .I(\current_shift_inst.phase_validZ0 ));
    Odrv12 I__5490 (
            .O(N__30164),
            .I(\current_shift_inst.phase_validZ0 ));
    Odrv4 I__5489 (
            .O(N__30161),
            .I(\current_shift_inst.phase_validZ0 ));
    InMux I__5488 (
            .O(N__30152),
            .I(N__30149));
    LocalMux I__5487 (
            .O(N__30149),
            .I(N__30146));
    Span4Mux_h I__5486 (
            .O(N__30146),
            .I(N__30143));
    Span4Mux_v I__5485 (
            .O(N__30143),
            .I(N__30140));
    Odrv4 I__5484 (
            .O(N__30140),
            .I(il_min_comp1_c));
    InMux I__5483 (
            .O(N__30137),
            .I(N__30134));
    LocalMux I__5482 (
            .O(N__30134),
            .I(il_min_comp1_D1));
    InMux I__5481 (
            .O(N__30131),
            .I(N__30128));
    LocalMux I__5480 (
            .O(N__30128),
            .I(il_min_comp2_D1));
    InMux I__5479 (
            .O(N__30125),
            .I(N__30121));
    InMux I__5478 (
            .O(N__30124),
            .I(N__30118));
    LocalMux I__5477 (
            .O(N__30121),
            .I(N__30113));
    LocalMux I__5476 (
            .O(N__30118),
            .I(N__30110));
    InMux I__5475 (
            .O(N__30117),
            .I(N__30105));
    InMux I__5474 (
            .O(N__30116),
            .I(N__30105));
    Span4Mux_h I__5473 (
            .O(N__30113),
            .I(N__30101));
    Span4Mux_v I__5472 (
            .O(N__30110),
            .I(N__30096));
    LocalMux I__5471 (
            .O(N__30105),
            .I(N__30096));
    InMux I__5470 (
            .O(N__30104),
            .I(N__30093));
    Odrv4 I__5469 (
            .O(N__30101),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_20 ));
    Odrv4 I__5468 (
            .O(N__30096),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_20 ));
    LocalMux I__5467 (
            .O(N__30093),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_20 ));
    CascadeMux I__5466 (
            .O(N__30086),
            .I(N__30083));
    InMux I__5465 (
            .O(N__30083),
            .I(N__30079));
    InMux I__5464 (
            .O(N__30082),
            .I(N__30076));
    LocalMux I__5463 (
            .O(N__30079),
            .I(N__30068));
    LocalMux I__5462 (
            .O(N__30076),
            .I(N__30068));
    InMux I__5461 (
            .O(N__30075),
            .I(N__30065));
    InMux I__5460 (
            .O(N__30074),
            .I(N__30060));
    InMux I__5459 (
            .O(N__30073),
            .I(N__30060));
    Span4Mux_v I__5458 (
            .O(N__30068),
            .I(N__30057));
    LocalMux I__5457 (
            .O(N__30065),
            .I(N__30054));
    LocalMux I__5456 (
            .O(N__30060),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    Odrv4 I__5455 (
            .O(N__30057),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    Odrv4 I__5454 (
            .O(N__30054),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    InMux I__5453 (
            .O(N__30047),
            .I(N__30044));
    LocalMux I__5452 (
            .O(N__30044),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__5451 (
            .O(N__30041),
            .I(N__30037));
    CascadeMux I__5450 (
            .O(N__30040),
            .I(N__30034));
    LocalMux I__5449 (
            .O(N__30037),
            .I(N__30031));
    InMux I__5448 (
            .O(N__30034),
            .I(N__30028));
    Span4Mux_v I__5447 (
            .O(N__30031),
            .I(N__30025));
    LocalMux I__5446 (
            .O(N__30028),
            .I(N__30021));
    Span4Mux_h I__5445 (
            .O(N__30025),
            .I(N__30018));
    InMux I__5444 (
            .O(N__30024),
            .I(N__30015));
    Odrv12 I__5443 (
            .O(N__30021),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__5442 (
            .O(N__30018),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__5441 (
            .O(N__30015),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    CascadeMux I__5440 (
            .O(N__30008),
            .I(N__30005));
    InMux I__5439 (
            .O(N__30005),
            .I(N__30002));
    LocalMux I__5438 (
            .O(N__30002),
            .I(N__29999));
    Span4Mux_h I__5437 (
            .O(N__29999),
            .I(N__29996));
    Odrv4 I__5436 (
            .O(N__29996),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__5435 (
            .O(N__29993),
            .I(N__29990));
    LocalMux I__5434 (
            .O(N__29990),
            .I(\current_shift_inst.un4_control_input_axb_17 ));
    InMux I__5433 (
            .O(N__29987),
            .I(N__29984));
    LocalMux I__5432 (
            .O(N__29984),
            .I(N__29981));
    Odrv4 I__5431 (
            .O(N__29981),
            .I(\current_shift_inst.un4_control_input_axb_21 ));
    InMux I__5430 (
            .O(N__29978),
            .I(N__29975));
    LocalMux I__5429 (
            .O(N__29975),
            .I(\current_shift_inst.un4_control_input_axb_26 ));
    InMux I__5428 (
            .O(N__29972),
            .I(N__29969));
    LocalMux I__5427 (
            .O(N__29969),
            .I(N__29965));
    InMux I__5426 (
            .O(N__29968),
            .I(N__29962));
    Span4Mux_v I__5425 (
            .O(N__29965),
            .I(N__29959));
    LocalMux I__5424 (
            .O(N__29962),
            .I(N__29956));
    Span4Mux_v I__5423 (
            .O(N__29959),
            .I(N__29953));
    Odrv4 I__5422 (
            .O(N__29956),
            .I(\current_shift_inst.z_31 ));
    Odrv4 I__5421 (
            .O(N__29953),
            .I(\current_shift_inst.z_31 ));
    CascadeMux I__5420 (
            .O(N__29948),
            .I(N__29944));
    InMux I__5419 (
            .O(N__29947),
            .I(N__29941));
    InMux I__5418 (
            .O(N__29944),
            .I(N__29938));
    LocalMux I__5417 (
            .O(N__29941),
            .I(N__29933));
    LocalMux I__5416 (
            .O(N__29938),
            .I(N__29933));
    Span4Mux_h I__5415 (
            .O(N__29933),
            .I(N__29930));
    Span4Mux_v I__5414 (
            .O(N__29930),
            .I(N__29927));
    Odrv4 I__5413 (
            .O(N__29927),
            .I(\current_shift_inst.z_i_31 ));
    InMux I__5412 (
            .O(N__29924),
            .I(N__29921));
    LocalMux I__5411 (
            .O(N__29921),
            .I(N__29918));
    Odrv4 I__5410 (
            .O(N__29918),
            .I(\current_shift_inst.un4_control_input_axb_30 ));
    InMux I__5409 (
            .O(N__29915),
            .I(N__29912));
    LocalMux I__5408 (
            .O(N__29912),
            .I(N__29909));
    Odrv4 I__5407 (
            .O(N__29909),
            .I(\current_shift_inst.un4_control_input_axb_27 ));
    InMux I__5406 (
            .O(N__29906),
            .I(N__29903));
    LocalMux I__5405 (
            .O(N__29903),
            .I(N__29900));
    Odrv4 I__5404 (
            .O(N__29900),
            .I(\current_shift_inst.un4_control_input_axb_29 ));
    InMux I__5403 (
            .O(N__29897),
            .I(N__29894));
    LocalMux I__5402 (
            .O(N__29894),
            .I(N__29891));
    Odrv4 I__5401 (
            .O(N__29891),
            .I(\current_shift_inst.un4_control_input_axb_28 ));
    InMux I__5400 (
            .O(N__29888),
            .I(N__29885));
    LocalMux I__5399 (
            .O(N__29885),
            .I(\current_shift_inst.un4_control_input_axb_12 ));
    InMux I__5398 (
            .O(N__29882),
            .I(N__29879));
    LocalMux I__5397 (
            .O(N__29879),
            .I(\current_shift_inst.un4_control_input_axb_16 ));
    InMux I__5396 (
            .O(N__29876),
            .I(N__29873));
    LocalMux I__5395 (
            .O(N__29873),
            .I(\current_shift_inst.un4_control_input_axb_20 ));
    InMux I__5394 (
            .O(N__29870),
            .I(N__29867));
    LocalMux I__5393 (
            .O(N__29867),
            .I(\current_shift_inst.un4_control_input_axb_18 ));
    InMux I__5392 (
            .O(N__29864),
            .I(N__29861));
    LocalMux I__5391 (
            .O(N__29861),
            .I(\current_shift_inst.un4_control_input_axb_23 ));
    InMux I__5390 (
            .O(N__29858),
            .I(N__29855));
    LocalMux I__5389 (
            .O(N__29855),
            .I(\current_shift_inst.un4_control_input_axb_19 ));
    InMux I__5388 (
            .O(N__29852),
            .I(N__29849));
    LocalMux I__5387 (
            .O(N__29849),
            .I(\current_shift_inst.un4_control_input_axb_25 ));
    InMux I__5386 (
            .O(N__29846),
            .I(N__29843));
    LocalMux I__5385 (
            .O(N__29843),
            .I(\current_shift_inst.un4_control_input_axb_22 ));
    InMux I__5384 (
            .O(N__29840),
            .I(N__29837));
    LocalMux I__5383 (
            .O(N__29837),
            .I(\current_shift_inst.un4_control_input_axb_24 ));
    InMux I__5382 (
            .O(N__29834),
            .I(N__29831));
    LocalMux I__5381 (
            .O(N__29831),
            .I(\current_shift_inst.un4_control_input_axb_4 ));
    InMux I__5380 (
            .O(N__29828),
            .I(N__29825));
    LocalMux I__5379 (
            .O(N__29825),
            .I(\current_shift_inst.un4_control_input_axb_5 ));
    InMux I__5378 (
            .O(N__29822),
            .I(N__29819));
    LocalMux I__5377 (
            .O(N__29819),
            .I(\current_shift_inst.un4_control_input_axb_6 ));
    CascadeMux I__5376 (
            .O(N__29816),
            .I(N__29813));
    InMux I__5375 (
            .O(N__29813),
            .I(N__29810));
    LocalMux I__5374 (
            .O(N__29810),
            .I(\current_shift_inst.un4_control_input_axb_7 ));
    CascadeMux I__5373 (
            .O(N__29807),
            .I(N__29804));
    InMux I__5372 (
            .O(N__29804),
            .I(N__29801));
    LocalMux I__5371 (
            .O(N__29801),
            .I(\current_shift_inst.un4_control_input_axb_8 ));
    InMux I__5370 (
            .O(N__29798),
            .I(N__29795));
    LocalMux I__5369 (
            .O(N__29795),
            .I(\current_shift_inst.un4_control_input_axb_13 ));
    InMux I__5368 (
            .O(N__29792),
            .I(N__29789));
    LocalMux I__5367 (
            .O(N__29789),
            .I(\current_shift_inst.un4_control_input_axb_15 ));
    InMux I__5366 (
            .O(N__29786),
            .I(N__29783));
    LocalMux I__5365 (
            .O(N__29783),
            .I(\current_shift_inst.un4_control_input_axb_9 ));
    InMux I__5364 (
            .O(N__29780),
            .I(N__29777));
    LocalMux I__5363 (
            .O(N__29777),
            .I(\current_shift_inst.un4_control_input_axb_10 ));
    InMux I__5362 (
            .O(N__29774),
            .I(N__29771));
    LocalMux I__5361 (
            .O(N__29771),
            .I(\current_shift_inst.un4_control_input_axb_11 ));
    InMux I__5360 (
            .O(N__29768),
            .I(N__29764));
    CascadeMux I__5359 (
            .O(N__29767),
            .I(N__29760));
    LocalMux I__5358 (
            .O(N__29764),
            .I(N__29757));
    InMux I__5357 (
            .O(N__29763),
            .I(N__29754));
    InMux I__5356 (
            .O(N__29760),
            .I(N__29751));
    Span4Mux_v I__5355 (
            .O(N__29757),
            .I(N__29748));
    LocalMux I__5354 (
            .O(N__29754),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    LocalMux I__5353 (
            .O(N__29751),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    Odrv4 I__5352 (
            .O(N__29748),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    InMux I__5351 (
            .O(N__29741),
            .I(N__29738));
    LocalMux I__5350 (
            .O(N__29738),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ));
    InMux I__5349 (
            .O(N__29735),
            .I(N__29732));
    LocalMux I__5348 (
            .O(N__29732),
            .I(\current_shift_inst.un4_control_input_axb_1 ));
    InMux I__5347 (
            .O(N__29729),
            .I(N__29726));
    LocalMux I__5346 (
            .O(N__29726),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ));
    InMux I__5345 (
            .O(N__29723),
            .I(N__29720));
    LocalMux I__5344 (
            .O(N__29720),
            .I(\current_shift_inst.un4_control_input_axb_2 ));
    InMux I__5343 (
            .O(N__29717),
            .I(N__29714));
    LocalMux I__5342 (
            .O(N__29714),
            .I(\current_shift_inst.un4_control_input_axb_14 ));
    InMux I__5341 (
            .O(N__29711),
            .I(N__29708));
    LocalMux I__5340 (
            .O(N__29708),
            .I(\current_shift_inst.un4_control_input_axb_3 ));
    CascadeMux I__5339 (
            .O(N__29705),
            .I(N__29701));
    CascadeMux I__5338 (
            .O(N__29704),
            .I(N__29698));
    InMux I__5337 (
            .O(N__29701),
            .I(N__29695));
    InMux I__5336 (
            .O(N__29698),
            .I(N__29690));
    LocalMux I__5335 (
            .O(N__29695),
            .I(N__29687));
    InMux I__5334 (
            .O(N__29694),
            .I(N__29684));
    InMux I__5333 (
            .O(N__29693),
            .I(N__29681));
    LocalMux I__5332 (
            .O(N__29690),
            .I(N__29678));
    Span4Mux_v I__5331 (
            .O(N__29687),
            .I(N__29675));
    LocalMux I__5330 (
            .O(N__29684),
            .I(N__29672));
    LocalMux I__5329 (
            .O(N__29681),
            .I(N__29669));
    Span4Mux_v I__5328 (
            .O(N__29678),
            .I(N__29666));
    Span4Mux_h I__5327 (
            .O(N__29675),
            .I(N__29659));
    Span4Mux_v I__5326 (
            .O(N__29672),
            .I(N__29659));
    Span4Mux_v I__5325 (
            .O(N__29669),
            .I(N__29659));
    Odrv4 I__5324 (
            .O(N__29666),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__5323 (
            .O(N__29659),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__5322 (
            .O(N__29654),
            .I(N__29651));
    InMux I__5321 (
            .O(N__29651),
            .I(N__29648));
    LocalMux I__5320 (
            .O(N__29648),
            .I(N__29645));
    Span4Mux_v I__5319 (
            .O(N__29645),
            .I(N__29642));
    Odrv4 I__5318 (
            .O(N__29642),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__5317 (
            .O(N__29639),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    InMux I__5316 (
            .O(N__29636),
            .I(N__29633));
    LocalMux I__5315 (
            .O(N__29633),
            .I(N__29628));
    InMux I__5314 (
            .O(N__29632),
            .I(N__29625));
    CascadeMux I__5313 (
            .O(N__29631),
            .I(N__29622));
    Span4Mux_v I__5312 (
            .O(N__29628),
            .I(N__29619));
    LocalMux I__5311 (
            .O(N__29625),
            .I(N__29616));
    InMux I__5310 (
            .O(N__29622),
            .I(N__29612));
    Span4Mux_h I__5309 (
            .O(N__29619),
            .I(N__29607));
    Span4Mux_h I__5308 (
            .O(N__29616),
            .I(N__29607));
    InMux I__5307 (
            .O(N__29615),
            .I(N__29604));
    LocalMux I__5306 (
            .O(N__29612),
            .I(N__29601));
    Odrv4 I__5305 (
            .O(N__29607),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__5304 (
            .O(N__29604),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv12 I__5303 (
            .O(N__29601),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__5302 (
            .O(N__29594),
            .I(N__29591));
    InMux I__5301 (
            .O(N__29591),
            .I(N__29588));
    LocalMux I__5300 (
            .O(N__29588),
            .I(N__29585));
    Sp12to4 I__5299 (
            .O(N__29585),
            .I(N__29582));
    Odrv12 I__5298 (
            .O(N__29582),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__5297 (
            .O(N__29579),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__5296 (
            .O(N__29576),
            .I(N__29572));
    CascadeMux I__5295 (
            .O(N__29575),
            .I(N__29569));
    InMux I__5294 (
            .O(N__29572),
            .I(N__29565));
    InMux I__5293 (
            .O(N__29569),
            .I(N__29562));
    CascadeMux I__5292 (
            .O(N__29568),
            .I(N__29558));
    LocalMux I__5291 (
            .O(N__29565),
            .I(N__29555));
    LocalMux I__5290 (
            .O(N__29562),
            .I(N__29552));
    InMux I__5289 (
            .O(N__29561),
            .I(N__29549));
    InMux I__5288 (
            .O(N__29558),
            .I(N__29546));
    Span4Mux_h I__5287 (
            .O(N__29555),
            .I(N__29543));
    Span4Mux_h I__5286 (
            .O(N__29552),
            .I(N__29538));
    LocalMux I__5285 (
            .O(N__29549),
            .I(N__29538));
    LocalMux I__5284 (
            .O(N__29546),
            .I(N__29535));
    Odrv4 I__5283 (
            .O(N__29543),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5282 (
            .O(N__29538),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5281 (
            .O(N__29535),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__5280 (
            .O(N__29528),
            .I(N__29525));
    InMux I__5279 (
            .O(N__29525),
            .I(N__29522));
    LocalMux I__5278 (
            .O(N__29522),
            .I(N__29519));
    Span4Mux_h I__5277 (
            .O(N__29519),
            .I(N__29516));
    Odrv4 I__5276 (
            .O(N__29516),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__5275 (
            .O(N__29513),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__5274 (
            .O(N__29510),
            .I(N__29503));
    CascadeMux I__5273 (
            .O(N__29509),
            .I(N__29500));
    CascadeMux I__5272 (
            .O(N__29508),
            .I(N__29496));
    CascadeMux I__5271 (
            .O(N__29507),
            .I(N__29492));
    CascadeMux I__5270 (
            .O(N__29506),
            .I(N__29488));
    LocalMux I__5269 (
            .O(N__29503),
            .I(N__29485));
    InMux I__5268 (
            .O(N__29500),
            .I(N__29470));
    InMux I__5267 (
            .O(N__29499),
            .I(N__29470));
    InMux I__5266 (
            .O(N__29496),
            .I(N__29470));
    InMux I__5265 (
            .O(N__29495),
            .I(N__29470));
    InMux I__5264 (
            .O(N__29492),
            .I(N__29470));
    InMux I__5263 (
            .O(N__29491),
            .I(N__29470));
    InMux I__5262 (
            .O(N__29488),
            .I(N__29470));
    Span4Mux_v I__5261 (
            .O(N__29485),
            .I(N__29467));
    LocalMux I__5260 (
            .O(N__29470),
            .I(N__29464));
    Span4Mux_v I__5259 (
            .O(N__29467),
            .I(N__29461));
    Span4Mux_h I__5258 (
            .O(N__29464),
            .I(N__29458));
    Odrv4 I__5257 (
            .O(N__29461),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    Odrv4 I__5256 (
            .O(N__29458),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    InMux I__5255 (
            .O(N__29453),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    CascadeMux I__5254 (
            .O(N__29450),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0_cascade_ ));
    InMux I__5253 (
            .O(N__29447),
            .I(N__29443));
    InMux I__5252 (
            .O(N__29446),
            .I(N__29440));
    LocalMux I__5251 (
            .O(N__29443),
            .I(N__29437));
    LocalMux I__5250 (
            .O(N__29440),
            .I(N__29434));
    Span4Mux_h I__5249 (
            .O(N__29437),
            .I(N__29431));
    Span4Mux_v I__5248 (
            .O(N__29434),
            .I(N__29428));
    Odrv4 I__5247 (
            .O(N__29431),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    Odrv4 I__5246 (
            .O(N__29428),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    InMux I__5245 (
            .O(N__29423),
            .I(N__29419));
    CascadeMux I__5244 (
            .O(N__29422),
            .I(N__29414));
    LocalMux I__5243 (
            .O(N__29419),
            .I(N__29411));
    InMux I__5242 (
            .O(N__29418),
            .I(N__29408));
    InMux I__5241 (
            .O(N__29417),
            .I(N__29405));
    InMux I__5240 (
            .O(N__29414),
            .I(N__29402));
    Span4Mux_h I__5239 (
            .O(N__29411),
            .I(N__29395));
    LocalMux I__5238 (
            .O(N__29408),
            .I(N__29395));
    LocalMux I__5237 (
            .O(N__29405),
            .I(N__29395));
    LocalMux I__5236 (
            .O(N__29402),
            .I(N__29392));
    Span4Mux_h I__5235 (
            .O(N__29395),
            .I(N__29389));
    Odrv12 I__5234 (
            .O(N__29392),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__5233 (
            .O(N__29389),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__5232 (
            .O(N__29384),
            .I(N__29381));
    InMux I__5231 (
            .O(N__29381),
            .I(N__29378));
    LocalMux I__5230 (
            .O(N__29378),
            .I(N__29375));
    Span4Mux_h I__5229 (
            .O(N__29375),
            .I(N__29372));
    Odrv4 I__5228 (
            .O(N__29372),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__5227 (
            .O(N__29369),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__5226 (
            .O(N__29366),
            .I(N__29363));
    InMux I__5225 (
            .O(N__29363),
            .I(N__29360));
    LocalMux I__5224 (
            .O(N__29360),
            .I(N__29357));
    Span4Mux_h I__5223 (
            .O(N__29357),
            .I(N__29351));
    InMux I__5222 (
            .O(N__29356),
            .I(N__29348));
    InMux I__5221 (
            .O(N__29355),
            .I(N__29343));
    InMux I__5220 (
            .O(N__29354),
            .I(N__29343));
    Odrv4 I__5219 (
            .O(N__29351),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__5218 (
            .O(N__29348),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__5217 (
            .O(N__29343),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    CascadeMux I__5216 (
            .O(N__29336),
            .I(N__29332));
    InMux I__5215 (
            .O(N__29335),
            .I(N__29329));
    InMux I__5214 (
            .O(N__29332),
            .I(N__29326));
    LocalMux I__5213 (
            .O(N__29329),
            .I(N__29323));
    LocalMux I__5212 (
            .O(N__29326),
            .I(N__29320));
    Span4Mux_v I__5211 (
            .O(N__29323),
            .I(N__29317));
    Span12Mux_v I__5210 (
            .O(N__29320),
            .I(N__29314));
    Odrv4 I__5209 (
            .O(N__29317),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    Odrv12 I__5208 (
            .O(N__29314),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    CascadeMux I__5207 (
            .O(N__29309),
            .I(N__29306));
    InMux I__5206 (
            .O(N__29306),
            .I(N__29303));
    LocalMux I__5205 (
            .O(N__29303),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__5204 (
            .O(N__29300),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__5203 (
            .O(N__29297),
            .I(N__29293));
    InMux I__5202 (
            .O(N__29296),
            .I(N__29288));
    InMux I__5201 (
            .O(N__29293),
            .I(N__29285));
    CascadeMux I__5200 (
            .O(N__29292),
            .I(N__29282));
    InMux I__5199 (
            .O(N__29291),
            .I(N__29279));
    LocalMux I__5198 (
            .O(N__29288),
            .I(N__29274));
    LocalMux I__5197 (
            .O(N__29285),
            .I(N__29274));
    InMux I__5196 (
            .O(N__29282),
            .I(N__29271));
    LocalMux I__5195 (
            .O(N__29279),
            .I(N__29268));
    Span4Mux_h I__5194 (
            .O(N__29274),
            .I(N__29265));
    LocalMux I__5193 (
            .O(N__29271),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5192 (
            .O(N__29268),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5191 (
            .O(N__29265),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__5190 (
            .O(N__29258),
            .I(N__29254));
    InMux I__5189 (
            .O(N__29257),
            .I(N__29251));
    InMux I__5188 (
            .O(N__29254),
            .I(N__29248));
    LocalMux I__5187 (
            .O(N__29251),
            .I(N__29245));
    LocalMux I__5186 (
            .O(N__29248),
            .I(N__29242));
    Span4Mux_h I__5185 (
            .O(N__29245),
            .I(N__29237));
    Span4Mux_h I__5184 (
            .O(N__29242),
            .I(N__29237));
    Odrv4 I__5183 (
            .O(N__29237),
            .I(\current_shift_inst.control_inputZ0Z_22 ));
    InMux I__5182 (
            .O(N__29234),
            .I(N__29231));
    LocalMux I__5181 (
            .O(N__29231),
            .I(N__29228));
    Odrv4 I__5180 (
            .O(N__29228),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__5179 (
            .O(N__29225),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__5178 (
            .O(N__29222),
            .I(N__29219));
    LocalMux I__5177 (
            .O(N__29219),
            .I(N__29213));
    InMux I__5176 (
            .O(N__29218),
            .I(N__29210));
    InMux I__5175 (
            .O(N__29217),
            .I(N__29207));
    InMux I__5174 (
            .O(N__29216),
            .I(N__29204));
    Span4Mux_h I__5173 (
            .O(N__29213),
            .I(N__29201));
    LocalMux I__5172 (
            .O(N__29210),
            .I(N__29198));
    LocalMux I__5171 (
            .O(N__29207),
            .I(N__29193));
    LocalMux I__5170 (
            .O(N__29204),
            .I(N__29193));
    Odrv4 I__5169 (
            .O(N__29201),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5168 (
            .O(N__29198),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5167 (
            .O(N__29193),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__5166 (
            .O(N__29186),
            .I(N__29182));
    InMux I__5165 (
            .O(N__29185),
            .I(N__29179));
    InMux I__5164 (
            .O(N__29182),
            .I(N__29176));
    LocalMux I__5163 (
            .O(N__29179),
            .I(N__29173));
    LocalMux I__5162 (
            .O(N__29176),
            .I(N__29170));
    Span4Mux_v I__5161 (
            .O(N__29173),
            .I(N__29165));
    Span4Mux_v I__5160 (
            .O(N__29170),
            .I(N__29165));
    Odrv4 I__5159 (
            .O(N__29165),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    CascadeMux I__5158 (
            .O(N__29162),
            .I(N__29159));
    InMux I__5157 (
            .O(N__29159),
            .I(N__29156));
    LocalMux I__5156 (
            .O(N__29156),
            .I(N__29153));
    Odrv4 I__5155 (
            .O(N__29153),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__5154 (
            .O(N__29150),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__5153 (
            .O(N__29147),
            .I(N__29143));
    InMux I__5152 (
            .O(N__29146),
            .I(N__29140));
    InMux I__5151 (
            .O(N__29143),
            .I(N__29137));
    LocalMux I__5150 (
            .O(N__29140),
            .I(N__29134));
    LocalMux I__5149 (
            .O(N__29137),
            .I(N__29131));
    Span12Mux_v I__5148 (
            .O(N__29134),
            .I(N__29128));
    Span4Mux_h I__5147 (
            .O(N__29131),
            .I(N__29125));
    Odrv12 I__5146 (
            .O(N__29128),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    Odrv4 I__5145 (
            .O(N__29125),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    InMux I__5144 (
            .O(N__29120),
            .I(bfn_11_13_0_));
    InMux I__5143 (
            .O(N__29117),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ));
    CascadeMux I__5142 (
            .O(N__29114),
            .I(N__29111));
    InMux I__5141 (
            .O(N__29111),
            .I(N__29108));
    LocalMux I__5140 (
            .O(N__29108),
            .I(N__29104));
    CascadeMux I__5139 (
            .O(N__29107),
            .I(N__29101));
    Span4Mux_v I__5138 (
            .O(N__29104),
            .I(N__29097));
    InMux I__5137 (
            .O(N__29101),
            .I(N__29094));
    CascadeMux I__5136 (
            .O(N__29100),
            .I(N__29090));
    Span4Mux_h I__5135 (
            .O(N__29097),
            .I(N__29087));
    LocalMux I__5134 (
            .O(N__29094),
            .I(N__29084));
    InMux I__5133 (
            .O(N__29093),
            .I(N__29079));
    InMux I__5132 (
            .O(N__29090),
            .I(N__29079));
    Odrv4 I__5131 (
            .O(N__29087),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__5130 (
            .O(N__29084),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__5129 (
            .O(N__29079),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__5128 (
            .O(N__29072),
            .I(N__29069));
    LocalMux I__5127 (
            .O(N__29069),
            .I(N__29066));
    Odrv4 I__5126 (
            .O(N__29066),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__5125 (
            .O(N__29063),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__5124 (
            .O(N__29060),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__5123 (
            .O(N__29057),
            .I(N__29053));
    InMux I__5122 (
            .O(N__29056),
            .I(N__29050));
    InMux I__5121 (
            .O(N__29053),
            .I(N__29047));
    LocalMux I__5120 (
            .O(N__29050),
            .I(N__29042));
    LocalMux I__5119 (
            .O(N__29047),
            .I(N__29039));
    InMux I__5118 (
            .O(N__29046),
            .I(N__29036));
    InMux I__5117 (
            .O(N__29045),
            .I(N__29033));
    Odrv12 I__5116 (
            .O(N__29042),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__5115 (
            .O(N__29039),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__5114 (
            .O(N__29036),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__5113 (
            .O(N__29033),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__5112 (
            .O(N__29024),
            .I(N__29020));
    InMux I__5111 (
            .O(N__29023),
            .I(N__29017));
    InMux I__5110 (
            .O(N__29020),
            .I(N__29014));
    LocalMux I__5109 (
            .O(N__29017),
            .I(N__29011));
    LocalMux I__5108 (
            .O(N__29014),
            .I(N__29008));
    Span4Mux_h I__5107 (
            .O(N__29011),
            .I(N__29005));
    Span12Mux_v I__5106 (
            .O(N__29008),
            .I(N__29002));
    Odrv4 I__5105 (
            .O(N__29005),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    Odrv12 I__5104 (
            .O(N__29002),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    CascadeMux I__5103 (
            .O(N__28997),
            .I(N__28994));
    InMux I__5102 (
            .O(N__28994),
            .I(N__28991));
    LocalMux I__5101 (
            .O(N__28991),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__5100 (
            .O(N__28988),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__5099 (
            .O(N__28985),
            .I(N__28981));
    InMux I__5098 (
            .O(N__28984),
            .I(N__28976));
    LocalMux I__5097 (
            .O(N__28981),
            .I(N__28973));
    InMux I__5096 (
            .O(N__28980),
            .I(N__28970));
    InMux I__5095 (
            .O(N__28979),
            .I(N__28967));
    LocalMux I__5094 (
            .O(N__28976),
            .I(N__28964));
    Odrv12 I__5093 (
            .O(N__28973),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__5092 (
            .O(N__28970),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__5091 (
            .O(N__28967),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__5090 (
            .O(N__28964),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__5089 (
            .O(N__28955),
            .I(N__28952));
    InMux I__5088 (
            .O(N__28952),
            .I(N__28948));
    InMux I__5087 (
            .O(N__28951),
            .I(N__28945));
    LocalMux I__5086 (
            .O(N__28948),
            .I(N__28942));
    LocalMux I__5085 (
            .O(N__28945),
            .I(N__28939));
    Span4Mux_h I__5084 (
            .O(N__28942),
            .I(N__28936));
    Span4Mux_v I__5083 (
            .O(N__28939),
            .I(N__28933));
    Span4Mux_h I__5082 (
            .O(N__28936),
            .I(N__28930));
    Odrv4 I__5081 (
            .O(N__28933),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    Odrv4 I__5080 (
            .O(N__28930),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    CascadeMux I__5079 (
            .O(N__28925),
            .I(N__28922));
    InMux I__5078 (
            .O(N__28922),
            .I(N__28919));
    LocalMux I__5077 (
            .O(N__28919),
            .I(N__28916));
    Odrv4 I__5076 (
            .O(N__28916),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__5075 (
            .O(N__28913),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__5074 (
            .O(N__28910),
            .I(N__28907));
    InMux I__5073 (
            .O(N__28907),
            .I(N__28903));
    InMux I__5072 (
            .O(N__28906),
            .I(N__28898));
    LocalMux I__5071 (
            .O(N__28903),
            .I(N__28895));
    InMux I__5070 (
            .O(N__28902),
            .I(N__28892));
    InMux I__5069 (
            .O(N__28901),
            .I(N__28889));
    LocalMux I__5068 (
            .O(N__28898),
            .I(N__28886));
    Odrv12 I__5067 (
            .O(N__28895),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__5066 (
            .O(N__28892),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__5065 (
            .O(N__28889),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__5064 (
            .O(N__28886),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__5063 (
            .O(N__28877),
            .I(N__28873));
    InMux I__5062 (
            .O(N__28876),
            .I(N__28870));
    InMux I__5061 (
            .O(N__28873),
            .I(N__28867));
    LocalMux I__5060 (
            .O(N__28870),
            .I(N__28864));
    LocalMux I__5059 (
            .O(N__28867),
            .I(N__28861));
    Span4Mux_h I__5058 (
            .O(N__28864),
            .I(N__28856));
    Span4Mux_h I__5057 (
            .O(N__28861),
            .I(N__28856));
    Span4Mux_h I__5056 (
            .O(N__28856),
            .I(N__28853));
    Odrv4 I__5055 (
            .O(N__28853),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    InMux I__5054 (
            .O(N__28850),
            .I(N__28847));
    LocalMux I__5053 (
            .O(N__28847),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__5052 (
            .O(N__28844),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__5051 (
            .O(N__28841),
            .I(N__28838));
    InMux I__5050 (
            .O(N__28838),
            .I(N__28834));
    CascadeMux I__5049 (
            .O(N__28837),
            .I(N__28830));
    LocalMux I__5048 (
            .O(N__28834),
            .I(N__28827));
    InMux I__5047 (
            .O(N__28833),
            .I(N__28823));
    InMux I__5046 (
            .O(N__28830),
            .I(N__28820));
    Span4Mux_h I__5045 (
            .O(N__28827),
            .I(N__28817));
    InMux I__5044 (
            .O(N__28826),
            .I(N__28814));
    LocalMux I__5043 (
            .O(N__28823),
            .I(N__28809));
    LocalMux I__5042 (
            .O(N__28820),
            .I(N__28809));
    Span4Mux_h I__5041 (
            .O(N__28817),
            .I(N__28806));
    LocalMux I__5040 (
            .O(N__28814),
            .I(N__28803));
    Span4Mux_h I__5039 (
            .O(N__28809),
            .I(N__28800));
    Odrv4 I__5038 (
            .O(N__28806),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv12 I__5037 (
            .O(N__28803),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__5036 (
            .O(N__28800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__5035 (
            .O(N__28793),
            .I(N__28789));
    InMux I__5034 (
            .O(N__28792),
            .I(N__28786));
    InMux I__5033 (
            .O(N__28789),
            .I(N__28783));
    LocalMux I__5032 (
            .O(N__28786),
            .I(N__28780));
    LocalMux I__5031 (
            .O(N__28783),
            .I(N__28777));
    Span4Mux_h I__5030 (
            .O(N__28780),
            .I(N__28774));
    Span4Mux_h I__5029 (
            .O(N__28777),
            .I(N__28771));
    Odrv4 I__5028 (
            .O(N__28774),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    Odrv4 I__5027 (
            .O(N__28771),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    CascadeMux I__5026 (
            .O(N__28766),
            .I(N__28763));
    InMux I__5025 (
            .O(N__28763),
            .I(N__28760));
    LocalMux I__5024 (
            .O(N__28760),
            .I(N__28757));
    Odrv4 I__5023 (
            .O(N__28757),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__5022 (
            .O(N__28754),
            .I(bfn_11_12_0_));
    InMux I__5021 (
            .O(N__28751),
            .I(N__28748));
    LocalMux I__5020 (
            .O(N__28748),
            .I(N__28744));
    InMux I__5019 (
            .O(N__28747),
            .I(N__28740));
    Span4Mux_v I__5018 (
            .O(N__28744),
            .I(N__28737));
    InMux I__5017 (
            .O(N__28743),
            .I(N__28733));
    LocalMux I__5016 (
            .O(N__28740),
            .I(N__28730));
    Span4Mux_h I__5015 (
            .O(N__28737),
            .I(N__28727));
    InMux I__5014 (
            .O(N__28736),
            .I(N__28724));
    LocalMux I__5013 (
            .O(N__28733),
            .I(N__28719));
    Span4Mux_v I__5012 (
            .O(N__28730),
            .I(N__28719));
    Odrv4 I__5011 (
            .O(N__28727),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__5010 (
            .O(N__28724),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__5009 (
            .O(N__28719),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CascadeMux I__5008 (
            .O(N__28712),
            .I(N__28709));
    InMux I__5007 (
            .O(N__28709),
            .I(N__28705));
    InMux I__5006 (
            .O(N__28708),
            .I(N__28702));
    LocalMux I__5005 (
            .O(N__28705),
            .I(N__28699));
    LocalMux I__5004 (
            .O(N__28702),
            .I(N__28696));
    Span4Mux_h I__5003 (
            .O(N__28699),
            .I(N__28693));
    Odrv4 I__5002 (
            .O(N__28696),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    Odrv4 I__5001 (
            .O(N__28693),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    CascadeMux I__5000 (
            .O(N__28688),
            .I(N__28685));
    InMux I__4999 (
            .O(N__28685),
            .I(N__28682));
    LocalMux I__4998 (
            .O(N__28682),
            .I(N__28679));
    Span4Mux_h I__4997 (
            .O(N__28679),
            .I(N__28676));
    Odrv4 I__4996 (
            .O(N__28676),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__4995 (
            .O(N__28673),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ));
    InMux I__4994 (
            .O(N__28670),
            .I(N__28667));
    LocalMux I__4993 (
            .O(N__28667),
            .I(N__28664));
    Span4Mux_h I__4992 (
            .O(N__28664),
            .I(N__28660));
    InMux I__4991 (
            .O(N__28663),
            .I(N__28656));
    Span4Mux_h I__4990 (
            .O(N__28660),
            .I(N__28652));
    InMux I__4989 (
            .O(N__28659),
            .I(N__28649));
    LocalMux I__4988 (
            .O(N__28656),
            .I(N__28646));
    InMux I__4987 (
            .O(N__28655),
            .I(N__28643));
    Odrv4 I__4986 (
            .O(N__28652),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__4985 (
            .O(N__28649),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__4984 (
            .O(N__28646),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__4983 (
            .O(N__28643),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__4982 (
            .O(N__28634),
            .I(N__28630));
    InMux I__4981 (
            .O(N__28633),
            .I(N__28627));
    InMux I__4980 (
            .O(N__28630),
            .I(N__28624));
    LocalMux I__4979 (
            .O(N__28627),
            .I(N__28621));
    LocalMux I__4978 (
            .O(N__28624),
            .I(N__28618));
    Span4Mux_h I__4977 (
            .O(N__28621),
            .I(N__28615));
    Span4Mux_h I__4976 (
            .O(N__28618),
            .I(N__28612));
    Odrv4 I__4975 (
            .O(N__28615),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    Odrv4 I__4974 (
            .O(N__28612),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    CascadeMux I__4973 (
            .O(N__28607),
            .I(N__28604));
    InMux I__4972 (
            .O(N__28604),
            .I(N__28601));
    LocalMux I__4971 (
            .O(N__28601),
            .I(N__28598));
    Odrv4 I__4970 (
            .O(N__28598),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__4969 (
            .O(N__28595),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    InMux I__4968 (
            .O(N__28592),
            .I(N__28587));
    InMux I__4967 (
            .O(N__28591),
            .I(N__28584));
    InMux I__4966 (
            .O(N__28590),
            .I(N__28580));
    LocalMux I__4965 (
            .O(N__28587),
            .I(N__28577));
    LocalMux I__4964 (
            .O(N__28584),
            .I(N__28574));
    InMux I__4963 (
            .O(N__28583),
            .I(N__28571));
    LocalMux I__4962 (
            .O(N__28580),
            .I(N__28568));
    Span4Mux_h I__4961 (
            .O(N__28577),
            .I(N__28563));
    Span4Mux_h I__4960 (
            .O(N__28574),
            .I(N__28563));
    LocalMux I__4959 (
            .O(N__28571),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__4958 (
            .O(N__28568),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__4957 (
            .O(N__28563),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__4956 (
            .O(N__28556),
            .I(N__28552));
    InMux I__4955 (
            .O(N__28555),
            .I(N__28549));
    InMux I__4954 (
            .O(N__28552),
            .I(N__28546));
    LocalMux I__4953 (
            .O(N__28549),
            .I(N__28543));
    LocalMux I__4952 (
            .O(N__28546),
            .I(N__28540));
    Span4Mux_v I__4951 (
            .O(N__28543),
            .I(N__28537));
    Span4Mux_h I__4950 (
            .O(N__28540),
            .I(N__28534));
    Odrv4 I__4949 (
            .O(N__28537),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    Odrv4 I__4948 (
            .O(N__28534),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    InMux I__4947 (
            .O(N__28529),
            .I(N__28526));
    LocalMux I__4946 (
            .O(N__28526),
            .I(N__28523));
    Odrv12 I__4945 (
            .O(N__28523),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__4944 (
            .O(N__28520),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__4943 (
            .O(N__28517),
            .I(N__28514));
    LocalMux I__4942 (
            .O(N__28514),
            .I(N__28511));
    Span4Mux_h I__4941 (
            .O(N__28511),
            .I(N__28506));
    InMux I__4940 (
            .O(N__28510),
            .I(N__28500));
    InMux I__4939 (
            .O(N__28509),
            .I(N__28500));
    Span4Mux_h I__4938 (
            .O(N__28506),
            .I(N__28497));
    InMux I__4937 (
            .O(N__28505),
            .I(N__28494));
    LocalMux I__4936 (
            .O(N__28500),
            .I(N__28491));
    Odrv4 I__4935 (
            .O(N__28497),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4934 (
            .O(N__28494),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4933 (
            .O(N__28491),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__4932 (
            .O(N__28484),
            .I(N__28480));
    InMux I__4931 (
            .O(N__28483),
            .I(N__28477));
    InMux I__4930 (
            .O(N__28480),
            .I(N__28474));
    LocalMux I__4929 (
            .O(N__28477),
            .I(N__28471));
    LocalMux I__4928 (
            .O(N__28474),
            .I(N__28468));
    Span12Mux_v I__4927 (
            .O(N__28471),
            .I(N__28465));
    Span4Mux_h I__4926 (
            .O(N__28468),
            .I(N__28462));
    Odrv12 I__4925 (
            .O(N__28465),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    Odrv4 I__4924 (
            .O(N__28462),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__4923 (
            .O(N__28457),
            .I(N__28454));
    LocalMux I__4922 (
            .O(N__28454),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__4921 (
            .O(N__28451),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__4920 (
            .O(N__28448),
            .I(N__28445));
    InMux I__4919 (
            .O(N__28445),
            .I(N__28442));
    LocalMux I__4918 (
            .O(N__28442),
            .I(N__28437));
    InMux I__4917 (
            .O(N__28441),
            .I(N__28434));
    InMux I__4916 (
            .O(N__28440),
            .I(N__28431));
    Span4Mux_v I__4915 (
            .O(N__28437),
            .I(N__28424));
    LocalMux I__4914 (
            .O(N__28434),
            .I(N__28424));
    LocalMux I__4913 (
            .O(N__28431),
            .I(N__28424));
    Span4Mux_h I__4912 (
            .O(N__28424),
            .I(N__28420));
    InMux I__4911 (
            .O(N__28423),
            .I(N__28417));
    Odrv4 I__4910 (
            .O(N__28420),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__4909 (
            .O(N__28417),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__4908 (
            .O(N__28412),
            .I(N__28408));
    CascadeMux I__4907 (
            .O(N__28411),
            .I(N__28405));
    LocalMux I__4906 (
            .O(N__28408),
            .I(N__28402));
    InMux I__4905 (
            .O(N__28405),
            .I(N__28399));
    Span4Mux_h I__4904 (
            .O(N__28402),
            .I(N__28396));
    LocalMux I__4903 (
            .O(N__28399),
            .I(N__28393));
    Span4Mux_v I__4902 (
            .O(N__28396),
            .I(N__28388));
    Span4Mux_v I__4901 (
            .O(N__28393),
            .I(N__28388));
    Odrv4 I__4900 (
            .O(N__28388),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    CascadeMux I__4899 (
            .O(N__28385),
            .I(N__28382));
    InMux I__4898 (
            .O(N__28382),
            .I(N__28379));
    LocalMux I__4897 (
            .O(N__28379),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__4896 (
            .O(N__28376),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    InMux I__4895 (
            .O(N__28373),
            .I(N__28370));
    LocalMux I__4894 (
            .O(N__28370),
            .I(N__28367));
    Span4Mux_h I__4893 (
            .O(N__28367),
            .I(N__28362));
    InMux I__4892 (
            .O(N__28366),
            .I(N__28356));
    InMux I__4891 (
            .O(N__28365),
            .I(N__28356));
    Span4Mux_h I__4890 (
            .O(N__28362),
            .I(N__28353));
    InMux I__4889 (
            .O(N__28361),
            .I(N__28350));
    LocalMux I__4888 (
            .O(N__28356),
            .I(N__28347));
    Odrv4 I__4887 (
            .O(N__28353),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__4886 (
            .O(N__28350),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__4885 (
            .O(N__28347),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__4884 (
            .O(N__28340),
            .I(N__28336));
    InMux I__4883 (
            .O(N__28339),
            .I(N__28333));
    InMux I__4882 (
            .O(N__28336),
            .I(N__28330));
    LocalMux I__4881 (
            .O(N__28333),
            .I(N__28327));
    LocalMux I__4880 (
            .O(N__28330),
            .I(N__28324));
    Span4Mux_h I__4879 (
            .O(N__28327),
            .I(N__28319));
    Span4Mux_h I__4878 (
            .O(N__28324),
            .I(N__28319));
    Odrv4 I__4877 (
            .O(N__28319),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__4876 (
            .O(N__28316),
            .I(N__28313));
    LocalMux I__4875 (
            .O(N__28313),
            .I(N__28310));
    Odrv4 I__4874 (
            .O(N__28310),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__4873 (
            .O(N__28307),
            .I(bfn_11_11_0_));
    CascadeMux I__4872 (
            .O(N__28304),
            .I(N__28300));
    InMux I__4871 (
            .O(N__28303),
            .I(N__28297));
    InMux I__4870 (
            .O(N__28300),
            .I(N__28293));
    LocalMux I__4869 (
            .O(N__28297),
            .I(N__28290));
    CascadeMux I__4868 (
            .O(N__28296),
            .I(N__28287));
    LocalMux I__4867 (
            .O(N__28293),
            .I(N__28281));
    Span4Mux_v I__4866 (
            .O(N__28290),
            .I(N__28281));
    InMux I__4865 (
            .O(N__28287),
            .I(N__28278));
    InMux I__4864 (
            .O(N__28286),
            .I(N__28275));
    Sp12to4 I__4863 (
            .O(N__28281),
            .I(N__28270));
    LocalMux I__4862 (
            .O(N__28278),
            .I(N__28270));
    LocalMux I__4861 (
            .O(N__28275),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__4860 (
            .O(N__28270),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__4859 (
            .O(N__28265),
            .I(N__28262));
    LocalMux I__4858 (
            .O(N__28262),
            .I(N__28258));
    CascadeMux I__4857 (
            .O(N__28261),
            .I(N__28255));
    Span4Mux_v I__4856 (
            .O(N__28258),
            .I(N__28252));
    InMux I__4855 (
            .O(N__28255),
            .I(N__28249));
    Span4Mux_v I__4854 (
            .O(N__28252),
            .I(N__28246));
    LocalMux I__4853 (
            .O(N__28249),
            .I(N__28243));
    Span4Mux_h I__4852 (
            .O(N__28246),
            .I(N__28240));
    Span4Mux_h I__4851 (
            .O(N__28243),
            .I(N__28237));
    Odrv4 I__4850 (
            .O(N__28240),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    Odrv4 I__4849 (
            .O(N__28237),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    CascadeMux I__4848 (
            .O(N__28232),
            .I(N__28229));
    InMux I__4847 (
            .O(N__28229),
            .I(N__28226));
    LocalMux I__4846 (
            .O(N__28226),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__4845 (
            .O(N__28223),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ));
    InMux I__4844 (
            .O(N__28220),
            .I(N__28216));
    CascadeMux I__4843 (
            .O(N__28219),
            .I(N__28213));
    LocalMux I__4842 (
            .O(N__28216),
            .I(N__28209));
    InMux I__4841 (
            .O(N__28213),
            .I(N__28206));
    InMux I__4840 (
            .O(N__28212),
            .I(N__28203));
    Span4Mux_h I__4839 (
            .O(N__28209),
            .I(N__28196));
    LocalMux I__4838 (
            .O(N__28206),
            .I(N__28196));
    LocalMux I__4837 (
            .O(N__28203),
            .I(N__28196));
    Span4Mux_h I__4836 (
            .O(N__28196),
            .I(N__28192));
    InMux I__4835 (
            .O(N__28195),
            .I(N__28189));
    Odrv4 I__4834 (
            .O(N__28192),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__4833 (
            .O(N__28189),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__4832 (
            .O(N__28184),
            .I(N__28180));
    CascadeMux I__4831 (
            .O(N__28183),
            .I(N__28177));
    LocalMux I__4830 (
            .O(N__28180),
            .I(N__28174));
    InMux I__4829 (
            .O(N__28177),
            .I(N__28171));
    Span4Mux_v I__4828 (
            .O(N__28174),
            .I(N__28168));
    LocalMux I__4827 (
            .O(N__28171),
            .I(N__28165));
    Span4Mux_h I__4826 (
            .O(N__28168),
            .I(N__28160));
    Span4Mux_h I__4825 (
            .O(N__28165),
            .I(N__28160));
    Odrv4 I__4824 (
            .O(N__28160),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    CascadeMux I__4823 (
            .O(N__28157),
            .I(N__28154));
    InMux I__4822 (
            .O(N__28154),
            .I(N__28151));
    LocalMux I__4821 (
            .O(N__28151),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__4820 (
            .O(N__28148),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    InMux I__4819 (
            .O(N__28145),
            .I(N__28141));
    InMux I__4818 (
            .O(N__28144),
            .I(N__28138));
    LocalMux I__4817 (
            .O(N__28141),
            .I(N__28135));
    LocalMux I__4816 (
            .O(N__28138),
            .I(N__28130));
    Span12Mux_s10_v I__4815 (
            .O(N__28135),
            .I(N__28127));
    InMux I__4814 (
            .O(N__28134),
            .I(N__28124));
    InMux I__4813 (
            .O(N__28133),
            .I(N__28121));
    Span4Mux_v I__4812 (
            .O(N__28130),
            .I(N__28118));
    Odrv12 I__4811 (
            .O(N__28127),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__4810 (
            .O(N__28124),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__4809 (
            .O(N__28121),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__4808 (
            .O(N__28118),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__4807 (
            .O(N__28109),
            .I(N__28105));
    InMux I__4806 (
            .O(N__28108),
            .I(N__28102));
    InMux I__4805 (
            .O(N__28105),
            .I(N__28099));
    LocalMux I__4804 (
            .O(N__28102),
            .I(N__28096));
    LocalMux I__4803 (
            .O(N__28099),
            .I(N__28093));
    Span4Mux_v I__4802 (
            .O(N__28096),
            .I(N__28090));
    Span4Mux_h I__4801 (
            .O(N__28093),
            .I(N__28087));
    Odrv4 I__4800 (
            .O(N__28090),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    Odrv4 I__4799 (
            .O(N__28087),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    CascadeMux I__4798 (
            .O(N__28082),
            .I(N__28079));
    InMux I__4797 (
            .O(N__28079),
            .I(N__28076));
    LocalMux I__4796 (
            .O(N__28076),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__4795 (
            .O(N__28073),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__4794 (
            .O(N__28070),
            .I(N__28066));
    CascadeMux I__4793 (
            .O(N__28069),
            .I(N__28063));
    LocalMux I__4792 (
            .O(N__28066),
            .I(N__28060));
    InMux I__4791 (
            .O(N__28063),
            .I(N__28057));
    Span4Mux_h I__4790 (
            .O(N__28060),
            .I(N__28051));
    LocalMux I__4789 (
            .O(N__28057),
            .I(N__28051));
    InMux I__4788 (
            .O(N__28056),
            .I(N__28047));
    Span4Mux_h I__4787 (
            .O(N__28051),
            .I(N__28044));
    InMux I__4786 (
            .O(N__28050),
            .I(N__28041));
    LocalMux I__4785 (
            .O(N__28047),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__4784 (
            .O(N__28044),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__4783 (
            .O(N__28041),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__4782 (
            .O(N__28034),
            .I(N__28031));
    InMux I__4781 (
            .O(N__28031),
            .I(N__28027));
    InMux I__4780 (
            .O(N__28030),
            .I(N__28024));
    LocalMux I__4779 (
            .O(N__28027),
            .I(N__28021));
    LocalMux I__4778 (
            .O(N__28024),
            .I(N__28018));
    Span4Mux_v I__4777 (
            .O(N__28021),
            .I(N__28015));
    Span4Mux_h I__4776 (
            .O(N__28018),
            .I(N__28012));
    Span4Mux_h I__4775 (
            .O(N__28015),
            .I(N__28009));
    Odrv4 I__4774 (
            .O(N__28012),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    Odrv4 I__4773 (
            .O(N__28009),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    InMux I__4772 (
            .O(N__28004),
            .I(N__28001));
    LocalMux I__4771 (
            .O(N__28001),
            .I(N__27998));
    Odrv4 I__4770 (
            .O(N__27998),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__4769 (
            .O(N__27995),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    InMux I__4768 (
            .O(N__27992),
            .I(N__27988));
    InMux I__4767 (
            .O(N__27991),
            .I(N__27985));
    LocalMux I__4766 (
            .O(N__27988),
            .I(N__27981));
    LocalMux I__4765 (
            .O(N__27985),
            .I(N__27978));
    InMux I__4764 (
            .O(N__27984),
            .I(N__27975));
    Span4Mux_v I__4763 (
            .O(N__27981),
            .I(N__27972));
    Odrv12 I__4762 (
            .O(N__27978),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__4761 (
            .O(N__27975),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__4760 (
            .O(N__27972),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__4759 (
            .O(N__27965),
            .I(N__27961));
    CascadeMux I__4758 (
            .O(N__27964),
            .I(N__27958));
    LocalMux I__4757 (
            .O(N__27961),
            .I(N__27955));
    InMux I__4756 (
            .O(N__27958),
            .I(N__27952));
    Span4Mux_v I__4755 (
            .O(N__27955),
            .I(N__27949));
    LocalMux I__4754 (
            .O(N__27952),
            .I(N__27946));
    Span4Mux_h I__4753 (
            .O(N__27949),
            .I(N__27941));
    Span4Mux_h I__4752 (
            .O(N__27946),
            .I(N__27941));
    Odrv4 I__4751 (
            .O(N__27941),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    CascadeMux I__4750 (
            .O(N__27938),
            .I(N__27935));
    InMux I__4749 (
            .O(N__27935),
            .I(N__27932));
    LocalMux I__4748 (
            .O(N__27932),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_axb_0 ));
    InMux I__4747 (
            .O(N__27929),
            .I(N__27926));
    LocalMux I__4746 (
            .O(N__27926),
            .I(N__27923));
    Span4Mux_h I__4745 (
            .O(N__27923),
            .I(N__27919));
    InMux I__4744 (
            .O(N__27922),
            .I(N__27915));
    Span4Mux_h I__4743 (
            .O(N__27919),
            .I(N__27912));
    InMux I__4742 (
            .O(N__27918),
            .I(N__27909));
    LocalMux I__4741 (
            .O(N__27915),
            .I(N__27906));
    Odrv4 I__4740 (
            .O(N__27912),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__4739 (
            .O(N__27909),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__4738 (
            .O(N__27906),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__4737 (
            .O(N__27899),
            .I(N__27896));
    InMux I__4736 (
            .O(N__27896),
            .I(N__27892));
    InMux I__4735 (
            .O(N__27895),
            .I(N__27889));
    LocalMux I__4734 (
            .O(N__27892),
            .I(N__27886));
    LocalMux I__4733 (
            .O(N__27889),
            .I(N__27883));
    Span4Mux_h I__4732 (
            .O(N__27886),
            .I(N__27880));
    Odrv4 I__4731 (
            .O(N__27883),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    Odrv4 I__4730 (
            .O(N__27880),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    CascadeMux I__4729 (
            .O(N__27875),
            .I(N__27872));
    InMux I__4728 (
            .O(N__27872),
            .I(N__27869));
    LocalMux I__4727 (
            .O(N__27869),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__4726 (
            .O(N__27866),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ));
    CascadeMux I__4725 (
            .O(N__27863),
            .I(N__27860));
    InMux I__4724 (
            .O(N__27860),
            .I(N__27856));
    InMux I__4723 (
            .O(N__27859),
            .I(N__27853));
    LocalMux I__4722 (
            .O(N__27856),
            .I(N__27850));
    LocalMux I__4721 (
            .O(N__27853),
            .I(N__27847));
    Span4Mux_h I__4720 (
            .O(N__27850),
            .I(N__27844));
    Odrv4 I__4719 (
            .O(N__27847),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    Odrv4 I__4718 (
            .O(N__27844),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__4717 (
            .O(N__27839),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__4716 (
            .O(N__27836),
            .I(N__27833));
    LocalMux I__4715 (
            .O(N__27833),
            .I(N__27829));
    InMux I__4714 (
            .O(N__27832),
            .I(N__27826));
    Span4Mux_v I__4713 (
            .O(N__27829),
            .I(N__27823));
    LocalMux I__4712 (
            .O(N__27826),
            .I(N__27820));
    Span4Mux_h I__4711 (
            .O(N__27823),
            .I(N__27817));
    Span4Mux_h I__4710 (
            .O(N__27820),
            .I(N__27814));
    Odrv4 I__4709 (
            .O(N__27817),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    Odrv4 I__4708 (
            .O(N__27814),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__4707 (
            .O(N__27809),
            .I(N__27806));
    LocalMux I__4706 (
            .O(N__27806),
            .I(N__27800));
    InMux I__4705 (
            .O(N__27805),
            .I(N__27797));
    InMux I__4704 (
            .O(N__27804),
            .I(N__27794));
    CascadeMux I__4703 (
            .O(N__27803),
            .I(N__27791));
    Span4Mux_v I__4702 (
            .O(N__27800),
            .I(N__27784));
    LocalMux I__4701 (
            .O(N__27797),
            .I(N__27784));
    LocalMux I__4700 (
            .O(N__27794),
            .I(N__27784));
    InMux I__4699 (
            .O(N__27791),
            .I(N__27781));
    Span4Mux_h I__4698 (
            .O(N__27784),
            .I(N__27778));
    LocalMux I__4697 (
            .O(N__27781),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__4696 (
            .O(N__27778),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__4695 (
            .O(N__27773),
            .I(N__27770));
    InMux I__4694 (
            .O(N__27770),
            .I(N__27767));
    LocalMux I__4693 (
            .O(N__27767),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__4692 (
            .O(N__27764),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    InMux I__4691 (
            .O(N__27761),
            .I(N__27755));
    InMux I__4690 (
            .O(N__27760),
            .I(N__27755));
    LocalMux I__4689 (
            .O(N__27755),
            .I(N__27751));
    InMux I__4688 (
            .O(N__27754),
            .I(N__27748));
    Span4Mux_v I__4687 (
            .O(N__27751),
            .I(N__27745));
    LocalMux I__4686 (
            .O(N__27748),
            .I(N__27741));
    Span4Mux_h I__4685 (
            .O(N__27745),
            .I(N__27738));
    InMux I__4684 (
            .O(N__27744),
            .I(N__27735));
    Odrv12 I__4683 (
            .O(N__27741),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__4682 (
            .O(N__27738),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__4681 (
            .O(N__27735),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__4680 (
            .O(N__27728),
            .I(N__27725));
    InMux I__4679 (
            .O(N__27725),
            .I(N__27722));
    LocalMux I__4678 (
            .O(N__27722),
            .I(N__27718));
    InMux I__4677 (
            .O(N__27721),
            .I(N__27715));
    Span4Mux_v I__4676 (
            .O(N__27718),
            .I(N__27712));
    LocalMux I__4675 (
            .O(N__27715),
            .I(N__27707));
    Span4Mux_h I__4674 (
            .O(N__27712),
            .I(N__27707));
    Odrv4 I__4673 (
            .O(N__27707),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    CascadeMux I__4672 (
            .O(N__27704),
            .I(N__27701));
    InMux I__4671 (
            .O(N__27701),
            .I(N__27698));
    LocalMux I__4670 (
            .O(N__27698),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__4669 (
            .O(N__27695),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__4668 (
            .O(N__27692),
            .I(N__27687));
    InMux I__4667 (
            .O(N__27691),
            .I(N__27684));
    InMux I__4666 (
            .O(N__27690),
            .I(N__27681));
    LocalMux I__4665 (
            .O(N__27687),
            .I(N__27678));
    LocalMux I__4664 (
            .O(N__27684),
            .I(N__27672));
    LocalMux I__4663 (
            .O(N__27681),
            .I(N__27672));
    Span4Mux_h I__4662 (
            .O(N__27678),
            .I(N__27669));
    InMux I__4661 (
            .O(N__27677),
            .I(N__27666));
    Span4Mux_h I__4660 (
            .O(N__27672),
            .I(N__27663));
    Odrv4 I__4659 (
            .O(N__27669),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__4658 (
            .O(N__27666),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__4657 (
            .O(N__27663),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__4656 (
            .O(N__27656),
            .I(N__27652));
    CascadeMux I__4655 (
            .O(N__27655),
            .I(N__27649));
    LocalMux I__4654 (
            .O(N__27652),
            .I(N__27646));
    InMux I__4653 (
            .O(N__27649),
            .I(N__27643));
    Span4Mux_h I__4652 (
            .O(N__27646),
            .I(N__27640));
    LocalMux I__4651 (
            .O(N__27643),
            .I(N__27637));
    Span4Mux_h I__4650 (
            .O(N__27640),
            .I(N__27634));
    Span12Mux_v I__4649 (
            .O(N__27637),
            .I(N__27631));
    Odrv4 I__4648 (
            .O(N__27634),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    Odrv12 I__4647 (
            .O(N__27631),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    CascadeMux I__4646 (
            .O(N__27626),
            .I(N__27623));
    InMux I__4645 (
            .O(N__27623),
            .I(N__27620));
    LocalMux I__4644 (
            .O(N__27620),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__4643 (
            .O(N__27617),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__4642 (
            .O(N__27614),
            .I(N__27609));
    CascadeMux I__4641 (
            .O(N__27613),
            .I(N__27606));
    CascadeMux I__4640 (
            .O(N__27612),
            .I(N__27603));
    InMux I__4639 (
            .O(N__27609),
            .I(N__27598));
    InMux I__4638 (
            .O(N__27606),
            .I(N__27595));
    InMux I__4637 (
            .O(N__27603),
            .I(N__27590));
    InMux I__4636 (
            .O(N__27602),
            .I(N__27590));
    InMux I__4635 (
            .O(N__27601),
            .I(N__27587));
    LocalMux I__4634 (
            .O(N__27598),
            .I(N__27584));
    LocalMux I__4633 (
            .O(N__27595),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__4632 (
            .O(N__27590),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__4631 (
            .O(N__27587),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv12 I__4630 (
            .O(N__27584),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__4629 (
            .O(N__27575),
            .I(N__27572));
    LocalMux I__4628 (
            .O(N__27572),
            .I(N__27569));
    Span4Mux_h I__4627 (
            .O(N__27569),
            .I(N__27564));
    InMux I__4626 (
            .O(N__27568),
            .I(N__27560));
    InMux I__4625 (
            .O(N__27567),
            .I(N__27557));
    Sp12to4 I__4624 (
            .O(N__27564),
            .I(N__27554));
    InMux I__4623 (
            .O(N__27563),
            .I(N__27551));
    LocalMux I__4622 (
            .O(N__27560),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__4621 (
            .O(N__27557),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__4620 (
            .O(N__27554),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__4619 (
            .O(N__27551),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__4618 (
            .O(N__27542),
            .I(N__27536));
    InMux I__4617 (
            .O(N__27541),
            .I(N__27533));
    InMux I__4616 (
            .O(N__27540),
            .I(N__27530));
    InMux I__4615 (
            .O(N__27539),
            .I(N__27527));
    LocalMux I__4614 (
            .O(N__27536),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__4613 (
            .O(N__27533),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__4612 (
            .O(N__27530),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__4611 (
            .O(N__27527),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    CEMux I__4610 (
            .O(N__27518),
            .I(N__27514));
    CEMux I__4609 (
            .O(N__27517),
            .I(N__27511));
    LocalMux I__4608 (
            .O(N__27514),
            .I(N__27508));
    LocalMux I__4607 (
            .O(N__27511),
            .I(N__27503));
    Span4Mux_v I__4606 (
            .O(N__27508),
            .I(N__27500));
    CEMux I__4605 (
            .O(N__27507),
            .I(N__27497));
    CEMux I__4604 (
            .O(N__27506),
            .I(N__27494));
    Span4Mux_v I__4603 (
            .O(N__27503),
            .I(N__27491));
    Span4Mux_h I__4602 (
            .O(N__27500),
            .I(N__27488));
    LocalMux I__4601 (
            .O(N__27497),
            .I(N__27485));
    LocalMux I__4600 (
            .O(N__27494),
            .I(N__27482));
    Odrv4 I__4599 (
            .O(N__27491),
            .I(\current_shift_inst.timer_s1.N_192_i ));
    Odrv4 I__4598 (
            .O(N__27488),
            .I(\current_shift_inst.timer_s1.N_192_i ));
    Odrv4 I__4597 (
            .O(N__27485),
            .I(\current_shift_inst.timer_s1.N_192_i ));
    Odrv12 I__4596 (
            .O(N__27482),
            .I(\current_shift_inst.timer_s1.N_192_i ));
    InMux I__4595 (
            .O(N__27473),
            .I(N__27467));
    InMux I__4594 (
            .O(N__27472),
            .I(N__27462));
    InMux I__4593 (
            .O(N__27471),
            .I(N__27462));
    InMux I__4592 (
            .O(N__27470),
            .I(N__27459));
    LocalMux I__4591 (
            .O(N__27467),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    LocalMux I__4590 (
            .O(N__27462),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    LocalMux I__4589 (
            .O(N__27459),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    InMux I__4588 (
            .O(N__27452),
            .I(N__27447));
    InMux I__4587 (
            .O(N__27451),
            .I(N__27443));
    InMux I__4586 (
            .O(N__27450),
            .I(N__27440));
    LocalMux I__4585 (
            .O(N__27447),
            .I(N__27437));
    InMux I__4584 (
            .O(N__27446),
            .I(N__27434));
    LocalMux I__4583 (
            .O(N__27443),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    LocalMux I__4582 (
            .O(N__27440),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv4 I__4581 (
            .O(N__27437),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    LocalMux I__4580 (
            .O(N__27434),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    IoInMux I__4579 (
            .O(N__27425),
            .I(N__27422));
    LocalMux I__4578 (
            .O(N__27422),
            .I(N__27419));
    IoSpan4Mux I__4577 (
            .O(N__27419),
            .I(N__27416));
    Span4Mux_s1_v I__4576 (
            .O(N__27416),
            .I(N__27413));
    Odrv4 I__4575 (
            .O(N__27413),
            .I(\current_shift_inst.timer_phase.N_188_i ));
    InMux I__4574 (
            .O(N__27410),
            .I(N__27407));
    LocalMux I__4573 (
            .O(N__27407),
            .I(N__27404));
    Span12Mux_h I__4572 (
            .O(N__27404),
            .I(N__27401));
    Odrv12 I__4571 (
            .O(N__27401),
            .I(il_max_comp2_c));
    InMux I__4570 (
            .O(N__27398),
            .I(N__27395));
    LocalMux I__4569 (
            .O(N__27395),
            .I(N__27392));
    Span4Mux_v I__4568 (
            .O(N__27392),
            .I(N__27389));
    Span4Mux_h I__4567 (
            .O(N__27389),
            .I(N__27386));
    Odrv4 I__4566 (
            .O(N__27386),
            .I(il_min_comp2_c));
    InMux I__4565 (
            .O(N__27383),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__4564 (
            .O(N__27380),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__4563 (
            .O(N__27377),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__4562 (
            .O(N__27374),
            .I(bfn_10_24_0_));
    InMux I__4561 (
            .O(N__27371),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__4560 (
            .O(N__27368),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__4559 (
            .O(N__27365),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__4558 (
            .O(N__27362),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__4557 (
            .O(N__27359),
            .I(N__27325));
    InMux I__4556 (
            .O(N__27358),
            .I(N__27325));
    InMux I__4555 (
            .O(N__27357),
            .I(N__27316));
    InMux I__4554 (
            .O(N__27356),
            .I(N__27316));
    InMux I__4553 (
            .O(N__27355),
            .I(N__27316));
    InMux I__4552 (
            .O(N__27354),
            .I(N__27316));
    InMux I__4551 (
            .O(N__27353),
            .I(N__27307));
    InMux I__4550 (
            .O(N__27352),
            .I(N__27307));
    InMux I__4549 (
            .O(N__27351),
            .I(N__27307));
    InMux I__4548 (
            .O(N__27350),
            .I(N__27307));
    InMux I__4547 (
            .O(N__27349),
            .I(N__27298));
    InMux I__4546 (
            .O(N__27348),
            .I(N__27298));
    InMux I__4545 (
            .O(N__27347),
            .I(N__27298));
    InMux I__4544 (
            .O(N__27346),
            .I(N__27298));
    InMux I__4543 (
            .O(N__27345),
            .I(N__27289));
    InMux I__4542 (
            .O(N__27344),
            .I(N__27289));
    InMux I__4541 (
            .O(N__27343),
            .I(N__27289));
    InMux I__4540 (
            .O(N__27342),
            .I(N__27289));
    InMux I__4539 (
            .O(N__27341),
            .I(N__27280));
    InMux I__4538 (
            .O(N__27340),
            .I(N__27280));
    InMux I__4537 (
            .O(N__27339),
            .I(N__27280));
    InMux I__4536 (
            .O(N__27338),
            .I(N__27280));
    InMux I__4535 (
            .O(N__27337),
            .I(N__27271));
    InMux I__4534 (
            .O(N__27336),
            .I(N__27271));
    InMux I__4533 (
            .O(N__27335),
            .I(N__27271));
    InMux I__4532 (
            .O(N__27334),
            .I(N__27271));
    InMux I__4531 (
            .O(N__27333),
            .I(N__27262));
    InMux I__4530 (
            .O(N__27332),
            .I(N__27262));
    InMux I__4529 (
            .O(N__27331),
            .I(N__27262));
    InMux I__4528 (
            .O(N__27330),
            .I(N__27262));
    LocalMux I__4527 (
            .O(N__27325),
            .I(N__27255));
    LocalMux I__4526 (
            .O(N__27316),
            .I(N__27255));
    LocalMux I__4525 (
            .O(N__27307),
            .I(N__27255));
    LocalMux I__4524 (
            .O(N__27298),
            .I(N__27242));
    LocalMux I__4523 (
            .O(N__27289),
            .I(N__27242));
    LocalMux I__4522 (
            .O(N__27280),
            .I(N__27242));
    LocalMux I__4521 (
            .O(N__27271),
            .I(N__27242));
    LocalMux I__4520 (
            .O(N__27262),
            .I(N__27242));
    Sp12to4 I__4519 (
            .O(N__27255),
            .I(N__27242));
    Odrv12 I__4518 (
            .O(N__27242),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__4517 (
            .O(N__27239),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__4516 (
            .O(N__27236),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__4515 (
            .O(N__27233),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__4514 (
            .O(N__27230),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__4513 (
            .O(N__27227),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__4512 (
            .O(N__27224),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__4511 (
            .O(N__27221),
            .I(bfn_10_23_0_));
    InMux I__4510 (
            .O(N__27218),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__4509 (
            .O(N__27215),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__4508 (
            .O(N__27212),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__4507 (
            .O(N__27209),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__4506 (
            .O(N__27206),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__4505 (
            .O(N__27203),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__4504 (
            .O(N__27200),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    InMux I__4503 (
            .O(N__27197),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__4502 (
            .O(N__27194),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__4501 (
            .O(N__27191),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__4500 (
            .O(N__27188),
            .I(bfn_10_22_0_));
    InMux I__4499 (
            .O(N__27185),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__4498 (
            .O(N__27182),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__4497 (
            .O(N__27179),
            .I(\current_shift_inst.un4_control_input_cry_26 ));
    InMux I__4496 (
            .O(N__27176),
            .I(\current_shift_inst.un4_control_input_cry_27 ));
    InMux I__4495 (
            .O(N__27173),
            .I(\current_shift_inst.un4_control_input_cry_28 ));
    InMux I__4494 (
            .O(N__27170),
            .I(N__27164));
    InMux I__4493 (
            .O(N__27169),
            .I(N__27164));
    LocalMux I__4492 (
            .O(N__27164),
            .I(N__27161));
    Span4Mux_h I__4491 (
            .O(N__27161),
            .I(N__27157));
    InMux I__4490 (
            .O(N__27160),
            .I(N__27154));
    Odrv4 I__4489 (
            .O(N__27157),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    LocalMux I__4488 (
            .O(N__27154),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    InMux I__4487 (
            .O(N__27149),
            .I(\current_shift_inst.un4_control_input_cry_29 ));
    CascadeMux I__4486 (
            .O(N__27146),
            .I(N__27143));
    InMux I__4485 (
            .O(N__27143),
            .I(N__27139));
    InMux I__4484 (
            .O(N__27142),
            .I(N__27136));
    LocalMux I__4483 (
            .O(N__27139),
            .I(N__27126));
    LocalMux I__4482 (
            .O(N__27136),
            .I(N__27126));
    InMux I__4481 (
            .O(N__27135),
            .I(N__27123));
    InMux I__4480 (
            .O(N__27134),
            .I(N__27120));
    InMux I__4479 (
            .O(N__27133),
            .I(N__27116));
    CascadeMux I__4478 (
            .O(N__27132),
            .I(N__27113));
    CascadeMux I__4477 (
            .O(N__27131),
            .I(N__27109));
    Span4Mux_v I__4476 (
            .O(N__27126),
            .I(N__27106));
    LocalMux I__4475 (
            .O(N__27123),
            .I(N__27103));
    LocalMux I__4474 (
            .O(N__27120),
            .I(N__27100));
    InMux I__4473 (
            .O(N__27119),
            .I(N__27097));
    LocalMux I__4472 (
            .O(N__27116),
            .I(N__27094));
    InMux I__4471 (
            .O(N__27113),
            .I(N__27087));
    InMux I__4470 (
            .O(N__27112),
            .I(N__27087));
    InMux I__4469 (
            .O(N__27109),
            .I(N__27087));
    Span4Mux_v I__4468 (
            .O(N__27106),
            .I(N__27082));
    Span4Mux_v I__4467 (
            .O(N__27103),
            .I(N__27082));
    Span4Mux_h I__4466 (
            .O(N__27100),
            .I(N__27079));
    LocalMux I__4465 (
            .O(N__27097),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__4464 (
            .O(N__27094),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__4463 (
            .O(N__27087),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__4462 (
            .O(N__27082),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__4461 (
            .O(N__27079),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__4460 (
            .O(N__27068),
            .I(\current_shift_inst.un4_control_input_cry_30 ));
    InMux I__4459 (
            .O(N__27065),
            .I(N__27059));
    InMux I__4458 (
            .O(N__27064),
            .I(N__27059));
    LocalMux I__4457 (
            .O(N__27059),
            .I(N__27056));
    Span4Mux_h I__4456 (
            .O(N__27056),
            .I(N__27052));
    InMux I__4455 (
            .O(N__27055),
            .I(N__27049));
    Odrv4 I__4454 (
            .O(N__27052),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    LocalMux I__4453 (
            .O(N__27049),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    InMux I__4452 (
            .O(N__27044),
            .I(N__27039));
    InMux I__4451 (
            .O(N__27043),
            .I(N__27033));
    InMux I__4450 (
            .O(N__27042),
            .I(N__27033));
    LocalMux I__4449 (
            .O(N__27039),
            .I(N__27030));
    InMux I__4448 (
            .O(N__27038),
            .I(N__27027));
    LocalMux I__4447 (
            .O(N__27033),
            .I(N__27024));
    Span4Mux_h I__4446 (
            .O(N__27030),
            .I(N__27021));
    LocalMux I__4445 (
            .O(N__27027),
            .I(N__27018));
    Odrv12 I__4444 (
            .O(N__27024),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    Odrv4 I__4443 (
            .O(N__27021),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    Odrv4 I__4442 (
            .O(N__27018),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    CascadeMux I__4441 (
            .O(N__27011),
            .I(N__27008));
    InMux I__4440 (
            .O(N__27008),
            .I(N__27002));
    InMux I__4439 (
            .O(N__27007),
            .I(N__27002));
    LocalMux I__4438 (
            .O(N__27002),
            .I(N__26997));
    CascadeMux I__4437 (
            .O(N__27001),
            .I(N__26994));
    InMux I__4436 (
            .O(N__27000),
            .I(N__26991));
    Span4Mux_h I__4435 (
            .O(N__26997),
            .I(N__26988));
    InMux I__4434 (
            .O(N__26994),
            .I(N__26985));
    LocalMux I__4433 (
            .O(N__26991),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    Odrv4 I__4432 (
            .O(N__26988),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    LocalMux I__4431 (
            .O(N__26985),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    InMux I__4430 (
            .O(N__26978),
            .I(N__26975));
    LocalMux I__4429 (
            .O(N__26975),
            .I(N__26972));
    Span4Mux_v I__4428 (
            .O(N__26972),
            .I(N__26969));
    Odrv4 I__4427 (
            .O(N__26969),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ));
    InMux I__4426 (
            .O(N__26966),
            .I(bfn_10_21_0_));
    InMux I__4425 (
            .O(N__26963),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__4424 (
            .O(N__26960),
            .I(N__26956));
    CascadeMux I__4423 (
            .O(N__26959),
            .I(N__26953));
    InMux I__4422 (
            .O(N__26956),
            .I(N__26948));
    InMux I__4421 (
            .O(N__26953),
            .I(N__26943));
    InMux I__4420 (
            .O(N__26952),
            .I(N__26943));
    CascadeMux I__4419 (
            .O(N__26951),
            .I(N__26940));
    LocalMux I__4418 (
            .O(N__26948),
            .I(N__26937));
    LocalMux I__4417 (
            .O(N__26943),
            .I(N__26934));
    InMux I__4416 (
            .O(N__26940),
            .I(N__26931));
    Odrv4 I__4415 (
            .O(N__26937),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    Odrv4 I__4414 (
            .O(N__26934),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    LocalMux I__4413 (
            .O(N__26931),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    InMux I__4412 (
            .O(N__26924),
            .I(\current_shift_inst.un4_control_input_cry_17 ));
    CascadeMux I__4411 (
            .O(N__26921),
            .I(N__26918));
    InMux I__4410 (
            .O(N__26918),
            .I(N__26915));
    LocalMux I__4409 (
            .O(N__26915),
            .I(N__26909));
    InMux I__4408 (
            .O(N__26914),
            .I(N__26904));
    InMux I__4407 (
            .O(N__26913),
            .I(N__26904));
    CascadeMux I__4406 (
            .O(N__26912),
            .I(N__26901));
    Span4Mux_v I__4405 (
            .O(N__26909),
            .I(N__26896));
    LocalMux I__4404 (
            .O(N__26904),
            .I(N__26896));
    InMux I__4403 (
            .O(N__26901),
            .I(N__26893));
    Odrv4 I__4402 (
            .O(N__26896),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    LocalMux I__4401 (
            .O(N__26893),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    InMux I__4400 (
            .O(N__26888),
            .I(\current_shift_inst.un4_control_input_cry_18 ));
    CascadeMux I__4399 (
            .O(N__26885),
            .I(N__26882));
    InMux I__4398 (
            .O(N__26882),
            .I(N__26879));
    LocalMux I__4397 (
            .O(N__26879),
            .I(N__26874));
    InMux I__4396 (
            .O(N__26878),
            .I(N__26869));
    InMux I__4395 (
            .O(N__26877),
            .I(N__26869));
    Span4Mux_v I__4394 (
            .O(N__26874),
            .I(N__26863));
    LocalMux I__4393 (
            .O(N__26869),
            .I(N__26863));
    CascadeMux I__4392 (
            .O(N__26868),
            .I(N__26860));
    Span4Mux_h I__4391 (
            .O(N__26863),
            .I(N__26857));
    InMux I__4390 (
            .O(N__26860),
            .I(N__26854));
    Odrv4 I__4389 (
            .O(N__26857),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    LocalMux I__4388 (
            .O(N__26854),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    InMux I__4387 (
            .O(N__26849),
            .I(\current_shift_inst.un4_control_input_cry_19 ));
    CascadeMux I__4386 (
            .O(N__26846),
            .I(N__26843));
    InMux I__4385 (
            .O(N__26843),
            .I(N__26837));
    InMux I__4384 (
            .O(N__26842),
            .I(N__26832));
    InMux I__4383 (
            .O(N__26841),
            .I(N__26832));
    CascadeMux I__4382 (
            .O(N__26840),
            .I(N__26829));
    LocalMux I__4381 (
            .O(N__26837),
            .I(N__26824));
    LocalMux I__4380 (
            .O(N__26832),
            .I(N__26824));
    InMux I__4379 (
            .O(N__26829),
            .I(N__26821));
    Odrv4 I__4378 (
            .O(N__26824),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    LocalMux I__4377 (
            .O(N__26821),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    InMux I__4376 (
            .O(N__26816),
            .I(\current_shift_inst.un4_control_input_cry_20 ));
    InMux I__4375 (
            .O(N__26813),
            .I(N__26807));
    InMux I__4374 (
            .O(N__26812),
            .I(N__26807));
    LocalMux I__4373 (
            .O(N__26807),
            .I(N__26803));
    InMux I__4372 (
            .O(N__26806),
            .I(N__26800));
    Span4Mux_h I__4371 (
            .O(N__26803),
            .I(N__26794));
    LocalMux I__4370 (
            .O(N__26800),
            .I(N__26794));
    InMux I__4369 (
            .O(N__26799),
            .I(N__26791));
    Odrv4 I__4368 (
            .O(N__26794),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    LocalMux I__4367 (
            .O(N__26791),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    InMux I__4366 (
            .O(N__26786),
            .I(\current_shift_inst.un4_control_input_cry_21 ));
    InMux I__4365 (
            .O(N__26783),
            .I(\current_shift_inst.un4_control_input_cry_22 ));
    InMux I__4364 (
            .O(N__26780),
            .I(\current_shift_inst.un4_control_input_cry_23 ));
    InMux I__4363 (
            .O(N__26777),
            .I(bfn_10_20_0_));
    InMux I__4362 (
            .O(N__26774),
            .I(\current_shift_inst.un4_control_input_cry_25 ));
    InMux I__4361 (
            .O(N__26771),
            .I(N__26766));
    InMux I__4360 (
            .O(N__26770),
            .I(N__26760));
    InMux I__4359 (
            .O(N__26769),
            .I(N__26760));
    LocalMux I__4358 (
            .O(N__26766),
            .I(N__26757));
    CascadeMux I__4357 (
            .O(N__26765),
            .I(N__26754));
    LocalMux I__4356 (
            .O(N__26760),
            .I(N__26751));
    Span4Mux_v I__4355 (
            .O(N__26757),
            .I(N__26748));
    InMux I__4354 (
            .O(N__26754),
            .I(N__26745));
    Odrv4 I__4353 (
            .O(N__26751),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    Odrv4 I__4352 (
            .O(N__26748),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    LocalMux I__4351 (
            .O(N__26745),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    InMux I__4350 (
            .O(N__26738),
            .I(bfn_10_18_0_));
    CascadeMux I__4349 (
            .O(N__26735),
            .I(N__26731));
    InMux I__4348 (
            .O(N__26734),
            .I(N__26727));
    InMux I__4347 (
            .O(N__26731),
            .I(N__26724));
    InMux I__4346 (
            .O(N__26730),
            .I(N__26721));
    LocalMux I__4345 (
            .O(N__26727),
            .I(N__26715));
    LocalMux I__4344 (
            .O(N__26724),
            .I(N__26715));
    LocalMux I__4343 (
            .O(N__26721),
            .I(N__26712));
    CascadeMux I__4342 (
            .O(N__26720),
            .I(N__26709));
    Span4Mux_v I__4341 (
            .O(N__26715),
            .I(N__26704));
    Span4Mux_v I__4340 (
            .O(N__26712),
            .I(N__26704));
    InMux I__4339 (
            .O(N__26709),
            .I(N__26701));
    Odrv4 I__4338 (
            .O(N__26704),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    LocalMux I__4337 (
            .O(N__26701),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    InMux I__4336 (
            .O(N__26696),
            .I(\current_shift_inst.un4_control_input_cry_9 ));
    CascadeMux I__4335 (
            .O(N__26693),
            .I(N__26690));
    InMux I__4334 (
            .O(N__26690),
            .I(N__26685));
    InMux I__4333 (
            .O(N__26689),
            .I(N__26682));
    InMux I__4332 (
            .O(N__26688),
            .I(N__26678));
    LocalMux I__4331 (
            .O(N__26685),
            .I(N__26673));
    LocalMux I__4330 (
            .O(N__26682),
            .I(N__26673));
    CascadeMux I__4329 (
            .O(N__26681),
            .I(N__26670));
    LocalMux I__4328 (
            .O(N__26678),
            .I(N__26665));
    Span4Mux_h I__4327 (
            .O(N__26673),
            .I(N__26665));
    InMux I__4326 (
            .O(N__26670),
            .I(N__26662));
    Odrv4 I__4325 (
            .O(N__26665),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    LocalMux I__4324 (
            .O(N__26662),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    InMux I__4323 (
            .O(N__26657),
            .I(\current_shift_inst.un4_control_input_cry_10 ));
    InMux I__4322 (
            .O(N__26654),
            .I(\current_shift_inst.un4_control_input_cry_11 ));
    InMux I__4321 (
            .O(N__26651),
            .I(\current_shift_inst.un4_control_input_cry_12 ));
    CascadeMux I__4320 (
            .O(N__26648),
            .I(N__26644));
    InMux I__4319 (
            .O(N__26647),
            .I(N__26640));
    InMux I__4318 (
            .O(N__26644),
            .I(N__26635));
    InMux I__4317 (
            .O(N__26643),
            .I(N__26635));
    LocalMux I__4316 (
            .O(N__26640),
            .I(N__26631));
    LocalMux I__4315 (
            .O(N__26635),
            .I(N__26628));
    CascadeMux I__4314 (
            .O(N__26634),
            .I(N__26625));
    Span4Mux_v I__4313 (
            .O(N__26631),
            .I(N__26622));
    Span4Mux_h I__4312 (
            .O(N__26628),
            .I(N__26619));
    InMux I__4311 (
            .O(N__26625),
            .I(N__26616));
    Odrv4 I__4310 (
            .O(N__26622),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    Odrv4 I__4309 (
            .O(N__26619),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    LocalMux I__4308 (
            .O(N__26616),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    InMux I__4307 (
            .O(N__26609),
            .I(\current_shift_inst.un4_control_input_cry_13 ));
    CascadeMux I__4306 (
            .O(N__26606),
            .I(N__26603));
    InMux I__4305 (
            .O(N__26603),
            .I(N__26600));
    LocalMux I__4304 (
            .O(N__26600),
            .I(N__26594));
    InMux I__4303 (
            .O(N__26599),
            .I(N__26591));
    InMux I__4302 (
            .O(N__26598),
            .I(N__26588));
    CascadeMux I__4301 (
            .O(N__26597),
            .I(N__26585));
    Sp12to4 I__4300 (
            .O(N__26594),
            .I(N__26578));
    LocalMux I__4299 (
            .O(N__26591),
            .I(N__26578));
    LocalMux I__4298 (
            .O(N__26588),
            .I(N__26578));
    InMux I__4297 (
            .O(N__26585),
            .I(N__26575));
    Odrv12 I__4296 (
            .O(N__26578),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    LocalMux I__4295 (
            .O(N__26575),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    InMux I__4294 (
            .O(N__26570),
            .I(\current_shift_inst.un4_control_input_cry_14 ));
    InMux I__4293 (
            .O(N__26567),
            .I(N__26562));
    InMux I__4292 (
            .O(N__26566),
            .I(N__26557));
    InMux I__4291 (
            .O(N__26565),
            .I(N__26557));
    LocalMux I__4290 (
            .O(N__26562),
            .I(N__26551));
    LocalMux I__4289 (
            .O(N__26557),
            .I(N__26551));
    InMux I__4288 (
            .O(N__26556),
            .I(N__26548));
    Odrv12 I__4287 (
            .O(N__26551),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    LocalMux I__4286 (
            .O(N__26548),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    InMux I__4285 (
            .O(N__26543),
            .I(\current_shift_inst.un4_control_input_cry_15 ));
    InMux I__4284 (
            .O(N__26540),
            .I(N__26535));
    InMux I__4283 (
            .O(N__26539),
            .I(N__26530));
    InMux I__4282 (
            .O(N__26538),
            .I(N__26530));
    LocalMux I__4281 (
            .O(N__26535),
            .I(N__26525));
    LocalMux I__4280 (
            .O(N__26530),
            .I(N__26525));
    Span4Mux_v I__4279 (
            .O(N__26525),
            .I(N__26521));
    InMux I__4278 (
            .O(N__26524),
            .I(N__26518));
    Odrv4 I__4277 (
            .O(N__26521),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    LocalMux I__4276 (
            .O(N__26518),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    InMux I__4275 (
            .O(N__26513),
            .I(bfn_10_19_0_));
    CascadeMux I__4274 (
            .O(N__26510),
            .I(N__26507));
    InMux I__4273 (
            .O(N__26507),
            .I(N__26504));
    LocalMux I__4272 (
            .O(N__26504),
            .I(N__26501));
    Span4Mux_h I__4271 (
            .O(N__26501),
            .I(N__26497));
    InMux I__4270 (
            .O(N__26500),
            .I(N__26494));
    Odrv4 I__4269 (
            .O(N__26497),
            .I(\current_shift_inst.un38_control_input_0 ));
    LocalMux I__4268 (
            .O(N__26494),
            .I(\current_shift_inst.un38_control_input_0 ));
    InMux I__4267 (
            .O(N__26489),
            .I(N__26485));
    InMux I__4266 (
            .O(N__26488),
            .I(N__26482));
    LocalMux I__4265 (
            .O(N__26485),
            .I(N__26479));
    LocalMux I__4264 (
            .O(N__26482),
            .I(N__26476));
    Span4Mux_v I__4263 (
            .O(N__26479),
            .I(N__26472));
    Span4Mux_h I__4262 (
            .O(N__26476),
            .I(N__26469));
    InMux I__4261 (
            .O(N__26475),
            .I(N__26466));
    Odrv4 I__4260 (
            .O(N__26472),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    Odrv4 I__4259 (
            .O(N__26469),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    LocalMux I__4258 (
            .O(N__26466),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    InMux I__4257 (
            .O(N__26459),
            .I(\current_shift_inst.un4_control_input_cry_1 ));
    CascadeMux I__4256 (
            .O(N__26456),
            .I(N__26452));
    InMux I__4255 (
            .O(N__26455),
            .I(N__26449));
    InMux I__4254 (
            .O(N__26452),
            .I(N__26445));
    LocalMux I__4253 (
            .O(N__26449),
            .I(N__26442));
    CascadeMux I__4252 (
            .O(N__26448),
            .I(N__26439));
    LocalMux I__4251 (
            .O(N__26445),
            .I(N__26436));
    Span4Mux_h I__4250 (
            .O(N__26442),
            .I(N__26433));
    InMux I__4249 (
            .O(N__26439),
            .I(N__26430));
    Odrv12 I__4248 (
            .O(N__26436),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    Odrv4 I__4247 (
            .O(N__26433),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    LocalMux I__4246 (
            .O(N__26430),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    InMux I__4245 (
            .O(N__26423),
            .I(\current_shift_inst.un4_control_input_cry_2 ));
    InMux I__4244 (
            .O(N__26420),
            .I(N__26417));
    LocalMux I__4243 (
            .O(N__26417),
            .I(N__26414));
    Span4Mux_h I__4242 (
            .O(N__26414),
            .I(N__26410));
    InMux I__4241 (
            .O(N__26413),
            .I(N__26407));
    Odrv4 I__4240 (
            .O(N__26410),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    LocalMux I__4239 (
            .O(N__26407),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    InMux I__4238 (
            .O(N__26402),
            .I(\current_shift_inst.un4_control_input_cry_3 ));
    InMux I__4237 (
            .O(N__26399),
            .I(N__26394));
    InMux I__4236 (
            .O(N__26398),
            .I(N__26389));
    InMux I__4235 (
            .O(N__26397),
            .I(N__26389));
    LocalMux I__4234 (
            .O(N__26394),
            .I(N__26383));
    LocalMux I__4233 (
            .O(N__26389),
            .I(N__26383));
    InMux I__4232 (
            .O(N__26388),
            .I(N__26380));
    Odrv12 I__4231 (
            .O(N__26383),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    LocalMux I__4230 (
            .O(N__26380),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    InMux I__4229 (
            .O(N__26375),
            .I(\current_shift_inst.un4_control_input_cry_4 ));
    CascadeMux I__4228 (
            .O(N__26372),
            .I(N__26369));
    InMux I__4227 (
            .O(N__26369),
            .I(N__26359));
    InMux I__4226 (
            .O(N__26368),
            .I(N__26359));
    InMux I__4225 (
            .O(N__26367),
            .I(N__26359));
    CascadeMux I__4224 (
            .O(N__26366),
            .I(N__26356));
    LocalMux I__4223 (
            .O(N__26359),
            .I(N__26353));
    InMux I__4222 (
            .O(N__26356),
            .I(N__26350));
    Odrv12 I__4221 (
            .O(N__26353),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    LocalMux I__4220 (
            .O(N__26350),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    InMux I__4219 (
            .O(N__26345),
            .I(\current_shift_inst.un4_control_input_cry_5 ));
    CascadeMux I__4218 (
            .O(N__26342),
            .I(N__26339));
    InMux I__4217 (
            .O(N__26339),
            .I(N__26331));
    InMux I__4216 (
            .O(N__26338),
            .I(N__26331));
    InMux I__4215 (
            .O(N__26337),
            .I(N__26328));
    CascadeMux I__4214 (
            .O(N__26336),
            .I(N__26325));
    LocalMux I__4213 (
            .O(N__26331),
            .I(N__26320));
    LocalMux I__4212 (
            .O(N__26328),
            .I(N__26320));
    InMux I__4211 (
            .O(N__26325),
            .I(N__26317));
    Odrv12 I__4210 (
            .O(N__26320),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    LocalMux I__4209 (
            .O(N__26317),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    InMux I__4208 (
            .O(N__26312),
            .I(\current_shift_inst.un4_control_input_cry_6 ));
    CascadeMux I__4207 (
            .O(N__26309),
            .I(N__26306));
    InMux I__4206 (
            .O(N__26306),
            .I(N__26300));
    InMux I__4205 (
            .O(N__26305),
            .I(N__26295));
    InMux I__4204 (
            .O(N__26304),
            .I(N__26295));
    CascadeMux I__4203 (
            .O(N__26303),
            .I(N__26292));
    LocalMux I__4202 (
            .O(N__26300),
            .I(N__26287));
    LocalMux I__4201 (
            .O(N__26295),
            .I(N__26287));
    InMux I__4200 (
            .O(N__26292),
            .I(N__26284));
    Odrv12 I__4199 (
            .O(N__26287),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    LocalMux I__4198 (
            .O(N__26284),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    InMux I__4197 (
            .O(N__26279),
            .I(\current_shift_inst.un4_control_input_cry_7 ));
    CascadeMux I__4196 (
            .O(N__26276),
            .I(N__26273));
    InMux I__4195 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__4194 (
            .O(N__26270),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ));
    CascadeMux I__4193 (
            .O(N__26267),
            .I(N__26264));
    InMux I__4192 (
            .O(N__26264),
            .I(N__26261));
    LocalMux I__4191 (
            .O(N__26261),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ));
    CascadeMux I__4190 (
            .O(N__26258),
            .I(N__26255));
    InMux I__4189 (
            .O(N__26255),
            .I(N__26252));
    LocalMux I__4188 (
            .O(N__26252),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ));
    CascadeMux I__4187 (
            .O(N__26249),
            .I(N__26246));
    InMux I__4186 (
            .O(N__26246),
            .I(N__26243));
    LocalMux I__4185 (
            .O(N__26243),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ));
    InMux I__4184 (
            .O(N__26240),
            .I(N__26236));
    CascadeMux I__4183 (
            .O(N__26239),
            .I(N__26233));
    LocalMux I__4182 (
            .O(N__26236),
            .I(N__26229));
    InMux I__4181 (
            .O(N__26233),
            .I(N__26224));
    InMux I__4180 (
            .O(N__26232),
            .I(N__26224));
    Span4Mux_v I__4179 (
            .O(N__26229),
            .I(N__26219));
    LocalMux I__4178 (
            .O(N__26224),
            .I(N__26219));
    Span4Mux_h I__4177 (
            .O(N__26219),
            .I(N__26215));
    InMux I__4176 (
            .O(N__26218),
            .I(N__26212));
    Span4Mux_v I__4175 (
            .O(N__26215),
            .I(N__26209));
    LocalMux I__4174 (
            .O(N__26212),
            .I(N__26206));
    Odrv4 I__4173 (
            .O(N__26209),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    Odrv4 I__4172 (
            .O(N__26206),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    InMux I__4171 (
            .O(N__26201),
            .I(N__26198));
    LocalMux I__4170 (
            .O(N__26198),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ));
    InMux I__4169 (
            .O(N__26195),
            .I(N__26189));
    InMux I__4168 (
            .O(N__26194),
            .I(N__26189));
    LocalMux I__4167 (
            .O(N__26189),
            .I(N__26184));
    InMux I__4166 (
            .O(N__26188),
            .I(N__26181));
    CascadeMux I__4165 (
            .O(N__26187),
            .I(N__26178));
    Span4Mux_h I__4164 (
            .O(N__26184),
            .I(N__26175));
    LocalMux I__4163 (
            .O(N__26181),
            .I(N__26172));
    InMux I__4162 (
            .O(N__26178),
            .I(N__26169));
    Span4Mux_v I__4161 (
            .O(N__26175),
            .I(N__26166));
    Span4Mux_h I__4160 (
            .O(N__26172),
            .I(N__26161));
    LocalMux I__4159 (
            .O(N__26169),
            .I(N__26161));
    Odrv4 I__4158 (
            .O(N__26166),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    Odrv4 I__4157 (
            .O(N__26161),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    InMux I__4156 (
            .O(N__26156),
            .I(N__26153));
    LocalMux I__4155 (
            .O(N__26153),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ));
    CascadeMux I__4154 (
            .O(N__26150),
            .I(N__26147));
    InMux I__4153 (
            .O(N__26147),
            .I(N__26141));
    InMux I__4152 (
            .O(N__26146),
            .I(N__26141));
    LocalMux I__4151 (
            .O(N__26141),
            .I(N__26136));
    InMux I__4150 (
            .O(N__26140),
            .I(N__26133));
    CascadeMux I__4149 (
            .O(N__26139),
            .I(N__26130));
    Span4Mux_h I__4148 (
            .O(N__26136),
            .I(N__26127));
    LocalMux I__4147 (
            .O(N__26133),
            .I(N__26124));
    InMux I__4146 (
            .O(N__26130),
            .I(N__26121));
    Span4Mux_v I__4145 (
            .O(N__26127),
            .I(N__26118));
    Span4Mux_h I__4144 (
            .O(N__26124),
            .I(N__26113));
    LocalMux I__4143 (
            .O(N__26121),
            .I(N__26113));
    Odrv4 I__4142 (
            .O(N__26118),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    Odrv4 I__4141 (
            .O(N__26113),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    InMux I__4140 (
            .O(N__26108),
            .I(N__26105));
    LocalMux I__4139 (
            .O(N__26105),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ));
    CascadeMux I__4138 (
            .O(N__26102),
            .I(N__26098));
    InMux I__4137 (
            .O(N__26101),
            .I(N__26090));
    InMux I__4136 (
            .O(N__26098),
            .I(N__26090));
    InMux I__4135 (
            .O(N__26097),
            .I(N__26090));
    LocalMux I__4134 (
            .O(N__26090),
            .I(N__26087));
    Span4Mux_v I__4133 (
            .O(N__26087),
            .I(N__26083));
    InMux I__4132 (
            .O(N__26086),
            .I(N__26080));
    Span4Mux_h I__4131 (
            .O(N__26083),
            .I(N__26077));
    LocalMux I__4130 (
            .O(N__26080),
            .I(N__26074));
    Odrv4 I__4129 (
            .O(N__26077),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    Odrv4 I__4128 (
            .O(N__26074),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    InMux I__4127 (
            .O(N__26069),
            .I(N__26062));
    InMux I__4126 (
            .O(N__26068),
            .I(N__26062));
    InMux I__4125 (
            .O(N__26067),
            .I(N__26059));
    LocalMux I__4124 (
            .O(N__26062),
            .I(N__26056));
    LocalMux I__4123 (
            .O(N__26059),
            .I(N__26053));
    Span4Mux_v I__4122 (
            .O(N__26056),
            .I(N__26050));
    Span4Mux_v I__4121 (
            .O(N__26053),
            .I(N__26044));
    Span4Mux_h I__4120 (
            .O(N__26050),
            .I(N__26044));
    InMux I__4119 (
            .O(N__26049),
            .I(N__26041));
    Span4Mux_h I__4118 (
            .O(N__26044),
            .I(N__26038));
    LocalMux I__4117 (
            .O(N__26041),
            .I(N__26035));
    Odrv4 I__4116 (
            .O(N__26038),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    Odrv4 I__4115 (
            .O(N__26035),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    InMux I__4114 (
            .O(N__26030),
            .I(N__26027));
    LocalMux I__4113 (
            .O(N__26027),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ));
    CascadeMux I__4112 (
            .O(N__26024),
            .I(N__26020));
    InMux I__4111 (
            .O(N__26023),
            .I(N__26012));
    InMux I__4110 (
            .O(N__26020),
            .I(N__26012));
    InMux I__4109 (
            .O(N__26019),
            .I(N__26012));
    LocalMux I__4108 (
            .O(N__26012),
            .I(N__26009));
    Span4Mux_h I__4107 (
            .O(N__26009),
            .I(N__26006));
    Span4Mux_v I__4106 (
            .O(N__26006),
            .I(N__26002));
    InMux I__4105 (
            .O(N__26005),
            .I(N__25999));
    Odrv4 I__4104 (
            .O(N__26002),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    LocalMux I__4103 (
            .O(N__25999),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    CascadeMux I__4102 (
            .O(N__25994),
            .I(N__25991));
    InMux I__4101 (
            .O(N__25991),
            .I(N__25984));
    InMux I__4100 (
            .O(N__25990),
            .I(N__25984));
    InMux I__4099 (
            .O(N__25989),
            .I(N__25981));
    LocalMux I__4098 (
            .O(N__25984),
            .I(N__25978));
    LocalMux I__4097 (
            .O(N__25981),
            .I(N__25975));
    Span4Mux_h I__4096 (
            .O(N__25978),
            .I(N__25972));
    Span12Mux_h I__4095 (
            .O(N__25975),
            .I(N__25968));
    Span4Mux_v I__4094 (
            .O(N__25972),
            .I(N__25965));
    InMux I__4093 (
            .O(N__25971),
            .I(N__25962));
    Odrv12 I__4092 (
            .O(N__25968),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    Odrv4 I__4091 (
            .O(N__25965),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    LocalMux I__4090 (
            .O(N__25962),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    InMux I__4089 (
            .O(N__25955),
            .I(N__25952));
    LocalMux I__4088 (
            .O(N__25952),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ));
    InMux I__4087 (
            .O(N__25949),
            .I(N__25946));
    LocalMux I__4086 (
            .O(N__25946),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ));
    CascadeMux I__4085 (
            .O(N__25943),
            .I(N__25940));
    InMux I__4084 (
            .O(N__25940),
            .I(N__25937));
    LocalMux I__4083 (
            .O(N__25937),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ));
    InMux I__4082 (
            .O(N__25934),
            .I(N__25929));
    InMux I__4081 (
            .O(N__25933),
            .I(N__25926));
    InMux I__4080 (
            .O(N__25932),
            .I(N__25923));
    LocalMux I__4079 (
            .O(N__25929),
            .I(N__25918));
    LocalMux I__4078 (
            .O(N__25926),
            .I(N__25918));
    LocalMux I__4077 (
            .O(N__25923),
            .I(N__25915));
    Span4Mux_v I__4076 (
            .O(N__25918),
            .I(N__25910));
    Span4Mux_h I__4075 (
            .O(N__25915),
            .I(N__25910));
    Span4Mux_v I__4074 (
            .O(N__25910),
            .I(N__25906));
    InMux I__4073 (
            .O(N__25909),
            .I(N__25903));
    Odrv4 I__4072 (
            .O(N__25906),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    LocalMux I__4071 (
            .O(N__25903),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    InMux I__4070 (
            .O(N__25898),
            .I(N__25895));
    LocalMux I__4069 (
            .O(N__25895),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ));
    InMux I__4068 (
            .O(N__25892),
            .I(N__25887));
    InMux I__4067 (
            .O(N__25891),
            .I(N__25884));
    InMux I__4066 (
            .O(N__25890),
            .I(N__25881));
    LocalMux I__4065 (
            .O(N__25887),
            .I(N__25877));
    LocalMux I__4064 (
            .O(N__25884),
            .I(N__25872));
    LocalMux I__4063 (
            .O(N__25881),
            .I(N__25872));
    CascadeMux I__4062 (
            .O(N__25880),
            .I(N__25869));
    Span4Mux_v I__4061 (
            .O(N__25877),
            .I(N__25866));
    Span4Mux_h I__4060 (
            .O(N__25872),
            .I(N__25863));
    InMux I__4059 (
            .O(N__25869),
            .I(N__25860));
    Span4Mux_h I__4058 (
            .O(N__25866),
            .I(N__25855));
    Span4Mux_v I__4057 (
            .O(N__25863),
            .I(N__25855));
    LocalMux I__4056 (
            .O(N__25860),
            .I(N__25852));
    Odrv4 I__4055 (
            .O(N__25855),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    Odrv4 I__4054 (
            .O(N__25852),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    InMux I__4053 (
            .O(N__25847),
            .I(N__25844));
    LocalMux I__4052 (
            .O(N__25844),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ));
    InMux I__4051 (
            .O(N__25841),
            .I(N__25838));
    LocalMux I__4050 (
            .O(N__25838),
            .I(N__25833));
    InMux I__4049 (
            .O(N__25837),
            .I(N__25830));
    InMux I__4048 (
            .O(N__25836),
            .I(N__25827));
    Span4Mux_v I__4047 (
            .O(N__25833),
            .I(N__25821));
    LocalMux I__4046 (
            .O(N__25830),
            .I(N__25821));
    LocalMux I__4045 (
            .O(N__25827),
            .I(N__25818));
    CascadeMux I__4044 (
            .O(N__25826),
            .I(N__25815));
    Span4Mux_h I__4043 (
            .O(N__25821),
            .I(N__25812));
    Span4Mux_h I__4042 (
            .O(N__25818),
            .I(N__25809));
    InMux I__4041 (
            .O(N__25815),
            .I(N__25806));
    Span4Mux_v I__4040 (
            .O(N__25812),
            .I(N__25803));
    Span4Mux_v I__4039 (
            .O(N__25809),
            .I(N__25798));
    LocalMux I__4038 (
            .O(N__25806),
            .I(N__25798));
    Odrv4 I__4037 (
            .O(N__25803),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    Odrv4 I__4036 (
            .O(N__25798),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    CascadeMux I__4035 (
            .O(N__25793),
            .I(N__25790));
    InMux I__4034 (
            .O(N__25790),
            .I(N__25787));
    LocalMux I__4033 (
            .O(N__25787),
            .I(N__25784));
    Odrv4 I__4032 (
            .O(N__25784),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ));
    CascadeMux I__4031 (
            .O(N__25781),
            .I(N__25778));
    InMux I__4030 (
            .O(N__25778),
            .I(N__25774));
    InMux I__4029 (
            .O(N__25777),
            .I(N__25771));
    LocalMux I__4028 (
            .O(N__25774),
            .I(N__25765));
    LocalMux I__4027 (
            .O(N__25771),
            .I(N__25765));
    InMux I__4026 (
            .O(N__25770),
            .I(N__25762));
    Span4Mux_v I__4025 (
            .O(N__25765),
            .I(N__25757));
    LocalMux I__4024 (
            .O(N__25762),
            .I(N__25757));
    Span4Mux_h I__4023 (
            .O(N__25757),
            .I(N__25754));
    Span4Mux_v I__4022 (
            .O(N__25754),
            .I(N__25750));
    InMux I__4021 (
            .O(N__25753),
            .I(N__25747));
    Odrv4 I__4020 (
            .O(N__25750),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    LocalMux I__4019 (
            .O(N__25747),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    InMux I__4018 (
            .O(N__25742),
            .I(N__25736));
    InMux I__4017 (
            .O(N__25741),
            .I(N__25731));
    InMux I__4016 (
            .O(N__25740),
            .I(N__25731));
    CascadeMux I__4015 (
            .O(N__25739),
            .I(N__25728));
    LocalMux I__4014 (
            .O(N__25736),
            .I(N__25725));
    LocalMux I__4013 (
            .O(N__25731),
            .I(N__25722));
    InMux I__4012 (
            .O(N__25728),
            .I(N__25719));
    Span12Mux_v I__4011 (
            .O(N__25725),
            .I(N__25716));
    Span4Mux_h I__4010 (
            .O(N__25722),
            .I(N__25711));
    LocalMux I__4009 (
            .O(N__25719),
            .I(N__25711));
    Odrv12 I__4008 (
            .O(N__25716),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    Odrv4 I__4007 (
            .O(N__25711),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    InMux I__4006 (
            .O(N__25706),
            .I(N__25703));
    LocalMux I__4005 (
            .O(N__25703),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ));
    InMux I__4004 (
            .O(N__25700),
            .I(N__25697));
    LocalMux I__4003 (
            .O(N__25697),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ));
    InMux I__4002 (
            .O(N__25694),
            .I(N__25691));
    LocalMux I__4001 (
            .O(N__25691),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ));
    CascadeMux I__4000 (
            .O(N__25688),
            .I(N__25685));
    InMux I__3999 (
            .O(N__25685),
            .I(N__25682));
    LocalMux I__3998 (
            .O(N__25682),
            .I(N__25677));
    InMux I__3997 (
            .O(N__25681),
            .I(N__25671));
    InMux I__3996 (
            .O(N__25680),
            .I(N__25671));
    Span4Mux_h I__3995 (
            .O(N__25677),
            .I(N__25668));
    InMux I__3994 (
            .O(N__25676),
            .I(N__25665));
    LocalMux I__3993 (
            .O(N__25671),
            .I(N__25662));
    Span4Mux_v I__3992 (
            .O(N__25668),
            .I(N__25657));
    LocalMux I__3991 (
            .O(N__25665),
            .I(N__25657));
    Odrv4 I__3990 (
            .O(N__25662),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    Odrv4 I__3989 (
            .O(N__25657),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    CascadeMux I__3988 (
            .O(N__25652),
            .I(N__25649));
    InMux I__3987 (
            .O(N__25649),
            .I(N__25646));
    LocalMux I__3986 (
            .O(N__25646),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ));
    InMux I__3985 (
            .O(N__25643),
            .I(N__25634));
    InMux I__3984 (
            .O(N__25642),
            .I(N__25634));
    InMux I__3983 (
            .O(N__25641),
            .I(N__25634));
    LocalMux I__3982 (
            .O(N__25634),
            .I(N__25631));
    Span4Mux_v I__3981 (
            .O(N__25631),
            .I(N__25627));
    InMux I__3980 (
            .O(N__25630),
            .I(N__25624));
    Span4Mux_h I__3979 (
            .O(N__25627),
            .I(N__25621));
    LocalMux I__3978 (
            .O(N__25624),
            .I(N__25618));
    Odrv4 I__3977 (
            .O(N__25621),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    Odrv4 I__3976 (
            .O(N__25618),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    CascadeMux I__3975 (
            .O(N__25613),
            .I(N__25609));
    CascadeMux I__3974 (
            .O(N__25612),
            .I(N__25606));
    InMux I__3973 (
            .O(N__25609),
            .I(N__25602));
    InMux I__3972 (
            .O(N__25606),
            .I(N__25597));
    InMux I__3971 (
            .O(N__25605),
            .I(N__25597));
    LocalMux I__3970 (
            .O(N__25602),
            .I(N__25594));
    LocalMux I__3969 (
            .O(N__25597),
            .I(N__25591));
    Span4Mux_v I__3968 (
            .O(N__25594),
            .I(N__25587));
    Span4Mux_h I__3967 (
            .O(N__25591),
            .I(N__25584));
    InMux I__3966 (
            .O(N__25590),
            .I(N__25581));
    Span4Mux_v I__3965 (
            .O(N__25587),
            .I(N__25578));
    Span4Mux_v I__3964 (
            .O(N__25584),
            .I(N__25573));
    LocalMux I__3963 (
            .O(N__25581),
            .I(N__25573));
    Odrv4 I__3962 (
            .O(N__25578),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    Odrv4 I__3961 (
            .O(N__25573),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    InMux I__3960 (
            .O(N__25568),
            .I(N__25565));
    LocalMux I__3959 (
            .O(N__25565),
            .I(N__25562));
    Odrv4 I__3958 (
            .O(N__25562),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ));
    CascadeMux I__3957 (
            .O(N__25559),
            .I(N__25556));
    InMux I__3956 (
            .O(N__25556),
            .I(N__25553));
    LocalMux I__3955 (
            .O(N__25553),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ));
    CascadeMux I__3954 (
            .O(N__25550),
            .I(N__25547));
    InMux I__3953 (
            .O(N__25547),
            .I(N__25544));
    LocalMux I__3952 (
            .O(N__25544),
            .I(N__25541));
    Odrv4 I__3951 (
            .O(N__25541),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ));
    CascadeMux I__3950 (
            .O(N__25538),
            .I(N__25535));
    InMux I__3949 (
            .O(N__25535),
            .I(N__25532));
    LocalMux I__3948 (
            .O(N__25532),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ));
    InMux I__3947 (
            .O(N__25529),
            .I(N__25526));
    LocalMux I__3946 (
            .O(N__25526),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ));
    CascadeMux I__3945 (
            .O(N__25523),
            .I(N__25520));
    InMux I__3944 (
            .O(N__25520),
            .I(N__25517));
    LocalMux I__3943 (
            .O(N__25517),
            .I(N__25514));
    Odrv4 I__3942 (
            .O(N__25514),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ));
    InMux I__3941 (
            .O(N__25511),
            .I(N__25508));
    LocalMux I__3940 (
            .O(N__25508),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ));
    InMux I__3939 (
            .O(N__25505),
            .I(N__25498));
    InMux I__3938 (
            .O(N__25504),
            .I(N__25498));
    InMux I__3937 (
            .O(N__25503),
            .I(N__25495));
    LocalMux I__3936 (
            .O(N__25498),
            .I(N__25492));
    LocalMux I__3935 (
            .O(N__25495),
            .I(N__25489));
    Span4Mux_v I__3934 (
            .O(N__25492),
            .I(N__25483));
    Span4Mux_v I__3933 (
            .O(N__25489),
            .I(N__25483));
    InMux I__3932 (
            .O(N__25488),
            .I(N__25480));
    Span4Mux_h I__3931 (
            .O(N__25483),
            .I(N__25477));
    LocalMux I__3930 (
            .O(N__25480),
            .I(N__25474));
    Odrv4 I__3929 (
            .O(N__25477),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    Odrv4 I__3928 (
            .O(N__25474),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    CascadeMux I__3927 (
            .O(N__25469),
            .I(N__25466));
    InMux I__3926 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__3925 (
            .O(N__25463),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ));
    InMux I__3924 (
            .O(N__25460),
            .I(N__25456));
    CascadeMux I__3923 (
            .O(N__25459),
            .I(N__25453));
    LocalMux I__3922 (
            .O(N__25456),
            .I(N__25450));
    InMux I__3921 (
            .O(N__25453),
            .I(N__25447));
    Span4Mux_v I__3920 (
            .O(N__25450),
            .I(N__25442));
    LocalMux I__3919 (
            .O(N__25447),
            .I(N__25442));
    Span4Mux_h I__3918 (
            .O(N__25442),
            .I(N__25439));
    Span4Mux_v I__3917 (
            .O(N__25439),
            .I(N__25436));
    Odrv4 I__3916 (
            .O(N__25436),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ));
    InMux I__3915 (
            .O(N__25433),
            .I(N__25430));
    LocalMux I__3914 (
            .O(N__25430),
            .I(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ));
    CascadeMux I__3913 (
            .O(N__25427),
            .I(N__25424));
    InMux I__3912 (
            .O(N__25424),
            .I(N__25421));
    LocalMux I__3911 (
            .O(N__25421),
            .I(N__25418));
    Odrv4 I__3910 (
            .O(N__25418),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ));
    InMux I__3909 (
            .O(N__25415),
            .I(N__25412));
    LocalMux I__3908 (
            .O(N__25412),
            .I(N__25409));
    Odrv4 I__3907 (
            .O(N__25409),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ));
    CascadeMux I__3906 (
            .O(N__25406),
            .I(N__25403));
    InMux I__3905 (
            .O(N__25403),
            .I(N__25400));
    LocalMux I__3904 (
            .O(N__25400),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ));
    CascadeMux I__3903 (
            .O(N__25397),
            .I(N__25394));
    InMux I__3902 (
            .O(N__25394),
            .I(N__25391));
    LocalMux I__3901 (
            .O(N__25391),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ));
    CascadeMux I__3900 (
            .O(N__25388),
            .I(N__25385));
    InMux I__3899 (
            .O(N__25385),
            .I(N__25382));
    LocalMux I__3898 (
            .O(N__25382),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ));
    CascadeMux I__3897 (
            .O(N__25379),
            .I(N__25376));
    InMux I__3896 (
            .O(N__25376),
            .I(N__25373));
    LocalMux I__3895 (
            .O(N__25373),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ));
    CascadeMux I__3894 (
            .O(N__25370),
            .I(N__25367));
    InMux I__3893 (
            .O(N__25367),
            .I(N__25364));
    LocalMux I__3892 (
            .O(N__25364),
            .I(N__25361));
    Odrv4 I__3891 (
            .O(N__25361),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ));
    InMux I__3890 (
            .O(N__25358),
            .I(N__25355));
    LocalMux I__3889 (
            .O(N__25355),
            .I(N__25352));
    Odrv4 I__3888 (
            .O(N__25352),
            .I(il_max_comp1_D1));
    CascadeMux I__3887 (
            .O(N__25349),
            .I(N__25346));
    InMux I__3886 (
            .O(N__25346),
            .I(N__25343));
    LocalMux I__3885 (
            .O(N__25343),
            .I(N__25340));
    Span4Mux_h I__3884 (
            .O(N__25340),
            .I(N__25337));
    Odrv4 I__3883 (
            .O(N__25337),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__3882 (
            .O(N__25334),
            .I(N__25331));
    InMux I__3881 (
            .O(N__25331),
            .I(N__25328));
    LocalMux I__3880 (
            .O(N__25328),
            .I(N__25325));
    Span4Mux_h I__3879 (
            .O(N__25325),
            .I(N__25322));
    Span4Mux_h I__3878 (
            .O(N__25322),
            .I(N__25319));
    Odrv4 I__3877 (
            .O(N__25319),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__3876 (
            .O(N__25316),
            .I(N__25313));
    InMux I__3875 (
            .O(N__25313),
            .I(N__25310));
    LocalMux I__3874 (
            .O(N__25310),
            .I(\current_shift_inst.z_5_30 ));
    InMux I__3873 (
            .O(N__25307),
            .I(N__25304));
    LocalMux I__3872 (
            .O(N__25304),
            .I(\current_shift_inst.z_5_cry_30_THRU_CO ));
    CascadeMux I__3871 (
            .O(N__25301),
            .I(N__25298));
    InMux I__3870 (
            .O(N__25298),
            .I(N__25294));
    InMux I__3869 (
            .O(N__25297),
            .I(N__25291));
    LocalMux I__3868 (
            .O(N__25294),
            .I(N__25288));
    LocalMux I__3867 (
            .O(N__25291),
            .I(N__25285));
    Span4Mux_h I__3866 (
            .O(N__25288),
            .I(N__25282));
    Odrv12 I__3865 (
            .O(N__25285),
            .I(\current_shift_inst.elapsed_time_ns_phase_31 ));
    Odrv4 I__3864 (
            .O(N__25282),
            .I(\current_shift_inst.elapsed_time_ns_phase_31 ));
    InMux I__3863 (
            .O(N__25277),
            .I(\current_shift_inst.z_cry_30 ));
    InMux I__3862 (
            .O(N__25274),
            .I(N__25271));
    LocalMux I__3861 (
            .O(N__25271),
            .I(N__25268));
    Odrv4 I__3860 (
            .O(N__25268),
            .I(\current_shift_inst.stop_timer_s1_RNOZ0Z_0 ));
    InMux I__3859 (
            .O(N__25265),
            .I(N__25260));
    InMux I__3858 (
            .O(N__25264),
            .I(N__25257));
    InMux I__3857 (
            .O(N__25263),
            .I(N__25254));
    LocalMux I__3856 (
            .O(N__25260),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    LocalMux I__3855 (
            .O(N__25257),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    LocalMux I__3854 (
            .O(N__25254),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    CascadeMux I__3853 (
            .O(N__25247),
            .I(N__25244));
    InMux I__3852 (
            .O(N__25244),
            .I(N__25241));
    LocalMux I__3851 (
            .O(N__25241),
            .I(\current_shift_inst.z_5_21 ));
    InMux I__3850 (
            .O(N__25238),
            .I(N__25235));
    LocalMux I__3849 (
            .O(N__25235),
            .I(\current_shift_inst.z_5_22 ));
    InMux I__3848 (
            .O(N__25232),
            .I(N__25229));
    LocalMux I__3847 (
            .O(N__25229),
            .I(\current_shift_inst.z_5_23 ));
    InMux I__3846 (
            .O(N__25226),
            .I(N__25223));
    LocalMux I__3845 (
            .O(N__25223),
            .I(N__25220));
    Odrv4 I__3844 (
            .O(N__25220),
            .I(\current_shift_inst.z_5_24 ));
    InMux I__3843 (
            .O(N__25217),
            .I(N__25214));
    LocalMux I__3842 (
            .O(N__25214),
            .I(\current_shift_inst.z_5_25 ));
    InMux I__3841 (
            .O(N__25211),
            .I(N__25208));
    LocalMux I__3840 (
            .O(N__25208),
            .I(\current_shift_inst.z_5_26 ));
    InMux I__3839 (
            .O(N__25205),
            .I(N__25202));
    LocalMux I__3838 (
            .O(N__25202),
            .I(\current_shift_inst.z_5_27 ));
    InMux I__3837 (
            .O(N__25199),
            .I(N__25196));
    LocalMux I__3836 (
            .O(N__25196),
            .I(\current_shift_inst.z_5_28 ));
    CascadeMux I__3835 (
            .O(N__25193),
            .I(N__25190));
    InMux I__3834 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__3833 (
            .O(N__25187),
            .I(\current_shift_inst.z_5_29 ));
    InMux I__3832 (
            .O(N__25184),
            .I(N__25181));
    LocalMux I__3831 (
            .O(N__25181),
            .I(\current_shift_inst.z_5_13 ));
    InMux I__3830 (
            .O(N__25178),
            .I(N__25175));
    LocalMux I__3829 (
            .O(N__25175),
            .I(\current_shift_inst.z_5_14 ));
    CascadeMux I__3828 (
            .O(N__25172),
            .I(N__25169));
    InMux I__3827 (
            .O(N__25169),
            .I(N__25166));
    LocalMux I__3826 (
            .O(N__25166),
            .I(\current_shift_inst.z_5_15 ));
    CascadeMux I__3825 (
            .O(N__25163),
            .I(N__25160));
    InMux I__3824 (
            .O(N__25160),
            .I(N__25157));
    LocalMux I__3823 (
            .O(N__25157),
            .I(N__25154));
    Span4Mux_v I__3822 (
            .O(N__25154),
            .I(N__25151));
    Odrv4 I__3821 (
            .O(N__25151),
            .I(\current_shift_inst.z_5_16 ));
    InMux I__3820 (
            .O(N__25148),
            .I(N__25145));
    LocalMux I__3819 (
            .O(N__25145),
            .I(\current_shift_inst.z_5_17 ));
    InMux I__3818 (
            .O(N__25142),
            .I(N__25139));
    LocalMux I__3817 (
            .O(N__25139),
            .I(\current_shift_inst.z_5_18 ));
    InMux I__3816 (
            .O(N__25136),
            .I(N__25133));
    LocalMux I__3815 (
            .O(N__25133),
            .I(\current_shift_inst.z_5_19 ));
    InMux I__3814 (
            .O(N__25130),
            .I(N__25127));
    LocalMux I__3813 (
            .O(N__25127),
            .I(\current_shift_inst.z_5_20 ));
    InMux I__3812 (
            .O(N__25124),
            .I(N__25121));
    LocalMux I__3811 (
            .O(N__25121),
            .I(\current_shift_inst.z_5_5 ));
    InMux I__3810 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__3809 (
            .O(N__25115),
            .I(\current_shift_inst.z_5_6 ));
    InMux I__3808 (
            .O(N__25112),
            .I(N__25109));
    LocalMux I__3807 (
            .O(N__25109),
            .I(\current_shift_inst.z_5_7 ));
    InMux I__3806 (
            .O(N__25106),
            .I(N__25103));
    LocalMux I__3805 (
            .O(N__25103),
            .I(N__25100));
    Odrv4 I__3804 (
            .O(N__25100),
            .I(\current_shift_inst.z_5_8 ));
    InMux I__3803 (
            .O(N__25097),
            .I(N__25094));
    LocalMux I__3802 (
            .O(N__25094),
            .I(\current_shift_inst.z_5_9 ));
    InMux I__3801 (
            .O(N__25091),
            .I(N__25088));
    LocalMux I__3800 (
            .O(N__25088),
            .I(\current_shift_inst.z_5_10 ));
    InMux I__3799 (
            .O(N__25085),
            .I(N__25082));
    LocalMux I__3798 (
            .O(N__25082),
            .I(\current_shift_inst.z_5_11 ));
    CascadeMux I__3797 (
            .O(N__25079),
            .I(N__25076));
    InMux I__3796 (
            .O(N__25076),
            .I(N__25073));
    LocalMux I__3795 (
            .O(N__25073),
            .I(\current_shift_inst.z_5_12 ));
    InMux I__3794 (
            .O(N__25070),
            .I(N__25067));
    LocalMux I__3793 (
            .O(N__25067),
            .I(N__25064));
    Odrv4 I__3792 (
            .O(N__25064),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ));
    CascadeMux I__3791 (
            .O(N__25061),
            .I(N__25058));
    InMux I__3790 (
            .O(N__25058),
            .I(N__25055));
    LocalMux I__3789 (
            .O(N__25055),
            .I(N__25052));
    Odrv4 I__3788 (
            .O(N__25052),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ));
    InMux I__3787 (
            .O(N__25049),
            .I(N__25046));
    LocalMux I__3786 (
            .O(N__25046),
            .I(\current_shift_inst.control_input_1_axb_23 ));
    InMux I__3785 (
            .O(N__25043),
            .I(\current_shift_inst.un38_control_input_0_cry_28 ));
    InMux I__3784 (
            .O(N__25040),
            .I(N__25037));
    LocalMux I__3783 (
            .O(N__25037),
            .I(N__25034));
    Span4Mux_v I__3782 (
            .O(N__25034),
            .I(N__25031));
    Odrv4 I__3781 (
            .O(N__25031),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ));
    CascadeMux I__3780 (
            .O(N__25028),
            .I(N__25024));
    InMux I__3779 (
            .O(N__25027),
            .I(N__25021));
    InMux I__3778 (
            .O(N__25024),
            .I(N__25018));
    LocalMux I__3777 (
            .O(N__25021),
            .I(N__25015));
    LocalMux I__3776 (
            .O(N__25018),
            .I(N__25012));
    Span4Mux_h I__3775 (
            .O(N__25015),
            .I(N__25009));
    Span4Mux_h I__3774 (
            .O(N__25012),
            .I(N__25006));
    Odrv4 I__3773 (
            .O(N__25009),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ));
    Odrv4 I__3772 (
            .O(N__25006),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ));
    InMux I__3771 (
            .O(N__25001),
            .I(N__24998));
    LocalMux I__3770 (
            .O(N__24998),
            .I(\current_shift_inst.control_input_1_axb_24 ));
    InMux I__3769 (
            .O(N__24995),
            .I(\current_shift_inst.un38_control_input_0_cry_29 ));
    InMux I__3768 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__3767 (
            .O(N__24989),
            .I(N__24986));
    Span4Mux_h I__3766 (
            .O(N__24986),
            .I(N__24983));
    Odrv4 I__3765 (
            .O(N__24983),
            .I(\current_shift_inst.un38_control_input_0_axb_31 ));
    CascadeMux I__3764 (
            .O(N__24980),
            .I(N__24977));
    InMux I__3763 (
            .O(N__24977),
            .I(N__24974));
    LocalMux I__3762 (
            .O(N__24974),
            .I(\current_shift_inst.control_input_1_cry_24_THRU_CO ));
    InMux I__3761 (
            .O(N__24971),
            .I(bfn_9_17_0_));
    CEMux I__3760 (
            .O(N__24968),
            .I(N__24963));
    CEMux I__3759 (
            .O(N__24967),
            .I(N__24960));
    CEMux I__3758 (
            .O(N__24966),
            .I(N__24956));
    LocalMux I__3757 (
            .O(N__24963),
            .I(N__24953));
    LocalMux I__3756 (
            .O(N__24960),
            .I(N__24949));
    CEMux I__3755 (
            .O(N__24959),
            .I(N__24946));
    LocalMux I__3754 (
            .O(N__24956),
            .I(N__24941));
    Span4Mux_v I__3753 (
            .O(N__24953),
            .I(N__24941));
    CEMux I__3752 (
            .O(N__24952),
            .I(N__24938));
    Span4Mux_v I__3751 (
            .O(N__24949),
            .I(N__24935));
    LocalMux I__3750 (
            .O(N__24946),
            .I(N__24928));
    Span4Mux_v I__3749 (
            .O(N__24941),
            .I(N__24928));
    LocalMux I__3748 (
            .O(N__24938),
            .I(N__24928));
    Odrv4 I__3747 (
            .O(N__24935),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    Odrv4 I__3746 (
            .O(N__24928),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    CascadeMux I__3745 (
            .O(N__24923),
            .I(N__24920));
    InMux I__3744 (
            .O(N__24920),
            .I(N__24917));
    LocalMux I__3743 (
            .O(N__24917),
            .I(G_406));
    InMux I__3742 (
            .O(N__24914),
            .I(N__24910));
    InMux I__3741 (
            .O(N__24913),
            .I(N__24904));
    LocalMux I__3740 (
            .O(N__24910),
            .I(N__24901));
    InMux I__3739 (
            .O(N__24909),
            .I(N__24897));
    InMux I__3738 (
            .O(N__24908),
            .I(N__24892));
    InMux I__3737 (
            .O(N__24907),
            .I(N__24892));
    LocalMux I__3736 (
            .O(N__24904),
            .I(N__24887));
    Span4Mux_h I__3735 (
            .O(N__24901),
            .I(N__24887));
    InMux I__3734 (
            .O(N__24900),
            .I(N__24884));
    LocalMux I__3733 (
            .O(N__24897),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    LocalMux I__3732 (
            .O(N__24892),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    Odrv4 I__3731 (
            .O(N__24887),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    LocalMux I__3730 (
            .O(N__24884),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    CascadeMux I__3729 (
            .O(N__24875),
            .I(N__24872));
    InMux I__3728 (
            .O(N__24872),
            .I(N__24869));
    LocalMux I__3727 (
            .O(N__24869),
            .I(G_405));
    InMux I__3726 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__3725 (
            .O(N__24863),
            .I(N__24860));
    Odrv4 I__3724 (
            .O(N__24860),
            .I(\current_shift_inst.z_5_2 ));
    CascadeMux I__3723 (
            .O(N__24857),
            .I(N__24854));
    InMux I__3722 (
            .O(N__24854),
            .I(N__24851));
    LocalMux I__3721 (
            .O(N__24851),
            .I(\current_shift_inst.z_5_3 ));
    CascadeMux I__3720 (
            .O(N__24848),
            .I(N__24845));
    InMux I__3719 (
            .O(N__24845),
            .I(N__24842));
    LocalMux I__3718 (
            .O(N__24842),
            .I(\current_shift_inst.z_5_4 ));
    InMux I__3717 (
            .O(N__24839),
            .I(N__24836));
    LocalMux I__3716 (
            .O(N__24836),
            .I(\current_shift_inst.control_input_1_axb_15 ));
    InMux I__3715 (
            .O(N__24833),
            .I(\current_shift_inst.un38_control_input_0_cry_20 ));
    InMux I__3714 (
            .O(N__24830),
            .I(N__24827));
    LocalMux I__3713 (
            .O(N__24827),
            .I(\current_shift_inst.control_input_1_axb_16 ));
    InMux I__3712 (
            .O(N__24824),
            .I(\current_shift_inst.un38_control_input_0_cry_21 ));
    InMux I__3711 (
            .O(N__24821),
            .I(N__24818));
    LocalMux I__3710 (
            .O(N__24818),
            .I(\current_shift_inst.control_input_1_axb_17 ));
    InMux I__3709 (
            .O(N__24815),
            .I(bfn_9_16_0_));
    InMux I__3708 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__3707 (
            .O(N__24809),
            .I(N__24806));
    Odrv4 I__3706 (
            .O(N__24806),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ));
    CascadeMux I__3705 (
            .O(N__24803),
            .I(N__24800));
    InMux I__3704 (
            .O(N__24800),
            .I(N__24797));
    LocalMux I__3703 (
            .O(N__24797),
            .I(N__24794));
    Odrv4 I__3702 (
            .O(N__24794),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ));
    InMux I__3701 (
            .O(N__24791),
            .I(N__24788));
    LocalMux I__3700 (
            .O(N__24788),
            .I(\current_shift_inst.control_input_1_axb_18 ));
    InMux I__3699 (
            .O(N__24785),
            .I(\current_shift_inst.un38_control_input_0_cry_23 ));
    InMux I__3698 (
            .O(N__24782),
            .I(N__24779));
    LocalMux I__3697 (
            .O(N__24779),
            .I(\current_shift_inst.control_input_1_axb_19 ));
    InMux I__3696 (
            .O(N__24776),
            .I(\current_shift_inst.un38_control_input_0_cry_24 ));
    InMux I__3695 (
            .O(N__24773),
            .I(N__24770));
    LocalMux I__3694 (
            .O(N__24770),
            .I(N__24767));
    Odrv4 I__3693 (
            .O(N__24767),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ));
    CascadeMux I__3692 (
            .O(N__24764),
            .I(N__24761));
    InMux I__3691 (
            .O(N__24761),
            .I(N__24758));
    LocalMux I__3690 (
            .O(N__24758),
            .I(N__24755));
    Odrv4 I__3689 (
            .O(N__24755),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ));
    InMux I__3688 (
            .O(N__24752),
            .I(N__24749));
    LocalMux I__3687 (
            .O(N__24749),
            .I(\current_shift_inst.control_input_1_axb_20 ));
    InMux I__3686 (
            .O(N__24746),
            .I(\current_shift_inst.un38_control_input_0_cry_25 ));
    InMux I__3685 (
            .O(N__24743),
            .I(N__24740));
    LocalMux I__3684 (
            .O(N__24740),
            .I(\current_shift_inst.control_input_1_axb_21 ));
    InMux I__3683 (
            .O(N__24737),
            .I(\current_shift_inst.un38_control_input_0_cry_26 ));
    CascadeMux I__3682 (
            .O(N__24734),
            .I(N__24731));
    InMux I__3681 (
            .O(N__24731),
            .I(N__24728));
    LocalMux I__3680 (
            .O(N__24728),
            .I(N__24725));
    Odrv4 I__3679 (
            .O(N__24725),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ));
    InMux I__3678 (
            .O(N__24722),
            .I(N__24719));
    LocalMux I__3677 (
            .O(N__24719),
            .I(\current_shift_inst.control_input_1_axb_22 ));
    InMux I__3676 (
            .O(N__24716),
            .I(\current_shift_inst.un38_control_input_0_cry_27 ));
    InMux I__3675 (
            .O(N__24713),
            .I(N__24710));
    LocalMux I__3674 (
            .O(N__24710),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__3673 (
            .O(N__24707),
            .I(\current_shift_inst.un38_control_input_0_cry_11 ));
    InMux I__3672 (
            .O(N__24704),
            .I(N__24701));
    LocalMux I__3671 (
            .O(N__24701),
            .I(N__24698));
    Span4Mux_h I__3670 (
            .O(N__24698),
            .I(N__24695));
    Odrv4 I__3669 (
            .O(N__24695),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ));
    InMux I__3668 (
            .O(N__24692),
            .I(N__24689));
    LocalMux I__3667 (
            .O(N__24689),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__3666 (
            .O(N__24686),
            .I(\current_shift_inst.un38_control_input_0_cry_12 ));
    InMux I__3665 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__3664 (
            .O(N__24680),
            .I(N__24677));
    Span4Mux_h I__3663 (
            .O(N__24677),
            .I(N__24674));
    Odrv4 I__3662 (
            .O(N__24674),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ));
    InMux I__3661 (
            .O(N__24671),
            .I(N__24668));
    LocalMux I__3660 (
            .O(N__24668),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__3659 (
            .O(N__24665),
            .I(\current_shift_inst.un38_control_input_0_cry_13 ));
    InMux I__3658 (
            .O(N__24662),
            .I(N__24659));
    LocalMux I__3657 (
            .O(N__24659),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__3656 (
            .O(N__24656),
            .I(bfn_9_15_0_));
    InMux I__3655 (
            .O(N__24653),
            .I(N__24650));
    LocalMux I__3654 (
            .O(N__24650),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__3653 (
            .O(N__24647),
            .I(\current_shift_inst.un38_control_input_0_cry_15 ));
    InMux I__3652 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__3651 (
            .O(N__24641),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__3650 (
            .O(N__24638),
            .I(\current_shift_inst.un38_control_input_0_cry_16 ));
    InMux I__3649 (
            .O(N__24635),
            .I(N__24632));
    LocalMux I__3648 (
            .O(N__24632),
            .I(\current_shift_inst.control_input_1_axb_12 ));
    InMux I__3647 (
            .O(N__24629),
            .I(\current_shift_inst.un38_control_input_0_cry_17 ));
    InMux I__3646 (
            .O(N__24626),
            .I(N__24623));
    LocalMux I__3645 (
            .O(N__24623),
            .I(\current_shift_inst.control_input_1_axb_13 ));
    InMux I__3644 (
            .O(N__24620),
            .I(\current_shift_inst.un38_control_input_0_cry_18 ));
    InMux I__3643 (
            .O(N__24617),
            .I(N__24614));
    LocalMux I__3642 (
            .O(N__24614),
            .I(\current_shift_inst.control_input_1_axb_14 ));
    InMux I__3641 (
            .O(N__24611),
            .I(\current_shift_inst.un38_control_input_0_cry_19 ));
    InMux I__3640 (
            .O(N__24608),
            .I(N__24605));
    LocalMux I__3639 (
            .O(N__24605),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__3638 (
            .O(N__24602),
            .I(\current_shift_inst.un38_control_input_0_cry_5 ));
    InMux I__3637 (
            .O(N__24599),
            .I(N__24596));
    LocalMux I__3636 (
            .O(N__24596),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__3635 (
            .O(N__24593),
            .I(bfn_9_14_0_));
    InMux I__3634 (
            .O(N__24590),
            .I(N__24587));
    LocalMux I__3633 (
            .O(N__24587),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__3632 (
            .O(N__24584),
            .I(\current_shift_inst.un38_control_input_0_cry_7 ));
    InMux I__3631 (
            .O(N__24581),
            .I(N__24578));
    LocalMux I__3630 (
            .O(N__24578),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__3629 (
            .O(N__24575),
            .I(\current_shift_inst.un38_control_input_0_cry_8 ));
    InMux I__3628 (
            .O(N__24572),
            .I(N__24569));
    LocalMux I__3627 (
            .O(N__24569),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__3626 (
            .O(N__24566),
            .I(\current_shift_inst.un38_control_input_0_cry_9 ));
    InMux I__3625 (
            .O(N__24563),
            .I(N__24560));
    LocalMux I__3624 (
            .O(N__24560),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__3623 (
            .O(N__24557),
            .I(\current_shift_inst.un38_control_input_0_cry_10 ));
    InMux I__3622 (
            .O(N__24554),
            .I(N__24551));
    LocalMux I__3621 (
            .O(N__24551),
            .I(\current_shift_inst.z_i_0_31 ));
    CascadeMux I__3620 (
            .O(N__24548),
            .I(N__24545));
    InMux I__3619 (
            .O(N__24545),
            .I(N__24542));
    LocalMux I__3618 (
            .O(N__24542),
            .I(N__24539));
    Span4Mux_v I__3617 (
            .O(N__24539),
            .I(N__24536));
    Odrv4 I__3616 (
            .O(N__24536),
            .I(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ));
    CascadeMux I__3615 (
            .O(N__24533),
            .I(N__24530));
    InMux I__3614 (
            .O(N__24530),
            .I(N__24527));
    LocalMux I__3613 (
            .O(N__24527),
            .I(N__24524));
    Span4Mux_h I__3612 (
            .O(N__24524),
            .I(N__24521));
    Odrv4 I__3611 (
            .O(N__24521),
            .I(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ));
    InMux I__3610 (
            .O(N__24518),
            .I(N__24515));
    LocalMux I__3609 (
            .O(N__24515),
            .I(N__24512));
    Span12Mux_v I__3608 (
            .O(N__24512),
            .I(N__24509));
    Odrv12 I__3607 (
            .O(N__24509),
            .I(\current_shift_inst.N_1620_i ));
    CascadeMux I__3606 (
            .O(N__24506),
            .I(N__24503));
    InMux I__3605 (
            .O(N__24503),
            .I(N__24500));
    LocalMux I__3604 (
            .O(N__24500),
            .I(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ));
    InMux I__3603 (
            .O(N__24497),
            .I(N__24494));
    LocalMux I__3602 (
            .O(N__24494),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    InMux I__3601 (
            .O(N__24491),
            .I(N__24486));
    InMux I__3600 (
            .O(N__24490),
            .I(N__24483));
    InMux I__3599 (
            .O(N__24489),
            .I(N__24480));
    LocalMux I__3598 (
            .O(N__24486),
            .I(N__24477));
    LocalMux I__3597 (
            .O(N__24483),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__3596 (
            .O(N__24480),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__3595 (
            .O(N__24477),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__3594 (
            .O(N__24470),
            .I(N__24465));
    InMux I__3593 (
            .O(N__24469),
            .I(N__24462));
    InMux I__3592 (
            .O(N__24468),
            .I(N__24459));
    LocalMux I__3591 (
            .O(N__24465),
            .I(N__24456));
    LocalMux I__3590 (
            .O(N__24462),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__3589 (
            .O(N__24459),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv12 I__3588 (
            .O(N__24456),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__3587 (
            .O(N__24449),
            .I(N__24446));
    LocalMux I__3586 (
            .O(N__24446),
            .I(\pwm_generator_inst.un1_counterlto2_0 ));
    CascadeMux I__3585 (
            .O(N__24443),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ));
    InMux I__3584 (
            .O(N__24440),
            .I(N__24437));
    LocalMux I__3583 (
            .O(N__24437),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    InMux I__3582 (
            .O(N__24434),
            .I(N__24431));
    LocalMux I__3581 (
            .O(N__24431),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__3580 (
            .O(N__24428),
            .I(N__24425));
    LocalMux I__3579 (
            .O(N__24425),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__3578 (
            .O(N__24422),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ));
    InMux I__3577 (
            .O(N__24419),
            .I(N__24416));
    LocalMux I__3576 (
            .O(N__24416),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__3575 (
            .O(N__24413),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__3574 (
            .O(N__24410),
            .I(N__24406));
    InMux I__3573 (
            .O(N__24409),
            .I(N__24402));
    LocalMux I__3572 (
            .O(N__24406),
            .I(N__24399));
    InMux I__3571 (
            .O(N__24405),
            .I(N__24396));
    LocalMux I__3570 (
            .O(N__24402),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__3569 (
            .O(N__24399),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__3568 (
            .O(N__24396),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__3567 (
            .O(N__24389),
            .I(N__24385));
    InMux I__3566 (
            .O(N__24388),
            .I(N__24381));
    LocalMux I__3565 (
            .O(N__24385),
            .I(N__24378));
    InMux I__3564 (
            .O(N__24384),
            .I(N__24375));
    LocalMux I__3563 (
            .O(N__24381),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__3562 (
            .O(N__24378),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__3561 (
            .O(N__24375),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__3560 (
            .O(N__24368),
            .I(N__24365));
    InMux I__3559 (
            .O(N__24365),
            .I(N__24361));
    InMux I__3558 (
            .O(N__24364),
            .I(N__24357));
    LocalMux I__3557 (
            .O(N__24361),
            .I(N__24354));
    InMux I__3556 (
            .O(N__24360),
            .I(N__24351));
    LocalMux I__3555 (
            .O(N__24357),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__3554 (
            .O(N__24354),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__3553 (
            .O(N__24351),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__3552 (
            .O(N__24344),
            .I(N__24341));
    LocalMux I__3551 (
            .O(N__24341),
            .I(N__24336));
    InMux I__3550 (
            .O(N__24340),
            .I(N__24333));
    InMux I__3549 (
            .O(N__24339),
            .I(N__24330));
    Odrv4 I__3548 (
            .O(N__24336),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__3547 (
            .O(N__24333),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__3546 (
            .O(N__24330),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__3545 (
            .O(N__24323),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__3544 (
            .O(N__24320),
            .I(N__24317));
    LocalMux I__3543 (
            .O(N__24317),
            .I(N__24312));
    InMux I__3542 (
            .O(N__24316),
            .I(N__24309));
    InMux I__3541 (
            .O(N__24315),
            .I(N__24306));
    Odrv4 I__3540 (
            .O(N__24312),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__3539 (
            .O(N__24309),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__3538 (
            .O(N__24306),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__3537 (
            .O(N__24299),
            .I(N__24281));
    InMux I__3536 (
            .O(N__24298),
            .I(N__24281));
    InMux I__3535 (
            .O(N__24297),
            .I(N__24281));
    InMux I__3534 (
            .O(N__24296),
            .I(N__24281));
    InMux I__3533 (
            .O(N__24295),
            .I(N__24272));
    InMux I__3532 (
            .O(N__24294),
            .I(N__24272));
    InMux I__3531 (
            .O(N__24293),
            .I(N__24272));
    InMux I__3530 (
            .O(N__24292),
            .I(N__24272));
    InMux I__3529 (
            .O(N__24291),
            .I(N__24267));
    InMux I__3528 (
            .O(N__24290),
            .I(N__24267));
    LocalMux I__3527 (
            .O(N__24281),
            .I(N__24262));
    LocalMux I__3526 (
            .O(N__24272),
            .I(N__24262));
    LocalMux I__3525 (
            .O(N__24267),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__3524 (
            .O(N__24262),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__3523 (
            .O(N__24257),
            .I(N__24252));
    InMux I__3522 (
            .O(N__24256),
            .I(N__24249));
    InMux I__3521 (
            .O(N__24255),
            .I(N__24246));
    LocalMux I__3520 (
            .O(N__24252),
            .I(N__24243));
    LocalMux I__3519 (
            .O(N__24249),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__3518 (
            .O(N__24246),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__3517 (
            .O(N__24243),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__3516 (
            .O(N__24236),
            .I(N__24231));
    InMux I__3515 (
            .O(N__24235),
            .I(N__24228));
    InMux I__3514 (
            .O(N__24234),
            .I(N__24225));
    LocalMux I__3513 (
            .O(N__24231),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__3512 (
            .O(N__24228),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__3511 (
            .O(N__24225),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__3510 (
            .O(N__24218),
            .I(N__24214));
    InMux I__3509 (
            .O(N__24217),
            .I(N__24210));
    LocalMux I__3508 (
            .O(N__24214),
            .I(N__24207));
    InMux I__3507 (
            .O(N__24213),
            .I(N__24204));
    LocalMux I__3506 (
            .O(N__24210),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__3505 (
            .O(N__24207),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__3504 (
            .O(N__24204),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__3503 (
            .O(N__24197),
            .I(N__24194));
    LocalMux I__3502 (
            .O(N__24194),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__3501 (
            .O(N__24191),
            .I(N__24188));
    LocalMux I__3500 (
            .O(N__24188),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    CascadeMux I__3499 (
            .O(N__24185),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ));
    InMux I__3498 (
            .O(N__24182),
            .I(N__24179));
    LocalMux I__3497 (
            .O(N__24179),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ));
    InMux I__3496 (
            .O(N__24176),
            .I(bfn_9_7_0_));
    InMux I__3495 (
            .O(N__24173),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__3494 (
            .O(N__24170),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__3493 (
            .O(N__24167),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__3492 (
            .O(N__24164),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__3491 (
            .O(N__24161),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__3490 (
            .O(N__24158),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__3489 (
            .O(N__24155),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__3488 (
            .O(N__24152),
            .I(bfn_9_8_0_));
    CascadeMux I__3487 (
            .O(N__24149),
            .I(N__24145));
    CascadeMux I__3486 (
            .O(N__24148),
            .I(N__24142));
    InMux I__3485 (
            .O(N__24145),
            .I(N__24139));
    InMux I__3484 (
            .O(N__24142),
            .I(N__24136));
    LocalMux I__3483 (
            .O(N__24139),
            .I(N__24132));
    LocalMux I__3482 (
            .O(N__24136),
            .I(N__24129));
    InMux I__3481 (
            .O(N__24135),
            .I(N__24126));
    Span4Mux_h I__3480 (
            .O(N__24132),
            .I(N__24123));
    Odrv4 I__3479 (
            .O(N__24129),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    LocalMux I__3478 (
            .O(N__24126),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    Odrv4 I__3477 (
            .O(N__24123),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    InMux I__3476 (
            .O(N__24116),
            .I(\current_shift_inst.timer_phase.counter_cry_24 ));
    CascadeMux I__3475 (
            .O(N__24113),
            .I(N__24109));
    InMux I__3474 (
            .O(N__24112),
            .I(N__24105));
    InMux I__3473 (
            .O(N__24109),
            .I(N__24102));
    InMux I__3472 (
            .O(N__24108),
            .I(N__24099));
    LocalMux I__3471 (
            .O(N__24105),
            .I(N__24094));
    LocalMux I__3470 (
            .O(N__24102),
            .I(N__24094));
    LocalMux I__3469 (
            .O(N__24099),
            .I(N__24089));
    Span4Mux_v I__3468 (
            .O(N__24094),
            .I(N__24089));
    Odrv4 I__3467 (
            .O(N__24089),
            .I(\current_shift_inst.timer_phase.counterZ0Z_26 ));
    InMux I__3466 (
            .O(N__24086),
            .I(\current_shift_inst.timer_phase.counter_cry_25 ));
    InMux I__3465 (
            .O(N__24083),
            .I(N__24076));
    InMux I__3464 (
            .O(N__24082),
            .I(N__24076));
    InMux I__3463 (
            .O(N__24081),
            .I(N__24073));
    LocalMux I__3462 (
            .O(N__24076),
            .I(N__24070));
    LocalMux I__3461 (
            .O(N__24073),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    Odrv4 I__3460 (
            .O(N__24070),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    InMux I__3459 (
            .O(N__24065),
            .I(\current_shift_inst.timer_phase.counter_cry_26 ));
    CascadeMux I__3458 (
            .O(N__24062),
            .I(N__24059));
    InMux I__3457 (
            .O(N__24059),
            .I(N__24055));
    InMux I__3456 (
            .O(N__24058),
            .I(N__24052));
    LocalMux I__3455 (
            .O(N__24055),
            .I(N__24049));
    LocalMux I__3454 (
            .O(N__24052),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    Odrv4 I__3453 (
            .O(N__24049),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    InMux I__3452 (
            .O(N__24044),
            .I(\current_shift_inst.timer_phase.counter_cry_27 ));
    InMux I__3451 (
            .O(N__24041),
            .I(\current_shift_inst.timer_phase.counter_cry_28 ));
    CascadeMux I__3450 (
            .O(N__24038),
            .I(N__24035));
    InMux I__3449 (
            .O(N__24035),
            .I(N__24031));
    InMux I__3448 (
            .O(N__24034),
            .I(N__24028));
    LocalMux I__3447 (
            .O(N__24031),
            .I(N__24025));
    LocalMux I__3446 (
            .O(N__24028),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    Odrv4 I__3445 (
            .O(N__24025),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    IoInMux I__3444 (
            .O(N__24020),
            .I(N__24017));
    LocalMux I__3443 (
            .O(N__24017),
            .I(N__24014));
    Span4Mux_s1_v I__3442 (
            .O(N__24014),
            .I(N__24011));
    Span4Mux_v I__3441 (
            .O(N__24011),
            .I(N__24008));
    Odrv4 I__3440 (
            .O(N__24008),
            .I(\current_shift_inst.timer_s1.N_187_i ));
    CEMux I__3439 (
            .O(N__24005),
            .I(N__24002));
    LocalMux I__3438 (
            .O(N__24002),
            .I(N__23997));
    CEMux I__3437 (
            .O(N__24001),
            .I(N__23994));
    CEMux I__3436 (
            .O(N__24000),
            .I(N__23991));
    Span4Mux_h I__3435 (
            .O(N__23997),
            .I(N__23986));
    LocalMux I__3434 (
            .O(N__23994),
            .I(N__23986));
    LocalMux I__3433 (
            .O(N__23991),
            .I(N__23982));
    Sp12to4 I__3432 (
            .O(N__23986),
            .I(N__23979));
    CEMux I__3431 (
            .O(N__23985),
            .I(N__23976));
    Odrv12 I__3430 (
            .O(N__23982),
            .I(\current_shift_inst.timer_phase.N_193_i ));
    Odrv12 I__3429 (
            .O(N__23979),
            .I(\current_shift_inst.timer_phase.N_193_i ));
    LocalMux I__3428 (
            .O(N__23976),
            .I(\current_shift_inst.timer_phase.N_193_i ));
    InMux I__3427 (
            .O(N__23969),
            .I(N__23931));
    InMux I__3426 (
            .O(N__23968),
            .I(N__23931));
    InMux I__3425 (
            .O(N__23967),
            .I(N__23931));
    InMux I__3424 (
            .O(N__23966),
            .I(N__23931));
    InMux I__3423 (
            .O(N__23965),
            .I(N__23922));
    InMux I__3422 (
            .O(N__23964),
            .I(N__23922));
    InMux I__3421 (
            .O(N__23963),
            .I(N__23922));
    InMux I__3420 (
            .O(N__23962),
            .I(N__23922));
    InMux I__3419 (
            .O(N__23961),
            .I(N__23913));
    InMux I__3418 (
            .O(N__23960),
            .I(N__23913));
    InMux I__3417 (
            .O(N__23959),
            .I(N__23913));
    InMux I__3416 (
            .O(N__23958),
            .I(N__23913));
    InMux I__3415 (
            .O(N__23957),
            .I(N__23904));
    InMux I__3414 (
            .O(N__23956),
            .I(N__23904));
    InMux I__3413 (
            .O(N__23955),
            .I(N__23904));
    InMux I__3412 (
            .O(N__23954),
            .I(N__23904));
    InMux I__3411 (
            .O(N__23953),
            .I(N__23895));
    InMux I__3410 (
            .O(N__23952),
            .I(N__23895));
    InMux I__3409 (
            .O(N__23951),
            .I(N__23895));
    InMux I__3408 (
            .O(N__23950),
            .I(N__23895));
    InMux I__3407 (
            .O(N__23949),
            .I(N__23886));
    InMux I__3406 (
            .O(N__23948),
            .I(N__23886));
    InMux I__3405 (
            .O(N__23947),
            .I(N__23886));
    InMux I__3404 (
            .O(N__23946),
            .I(N__23886));
    InMux I__3403 (
            .O(N__23945),
            .I(N__23881));
    InMux I__3402 (
            .O(N__23944),
            .I(N__23881));
    InMux I__3401 (
            .O(N__23943),
            .I(N__23872));
    InMux I__3400 (
            .O(N__23942),
            .I(N__23872));
    InMux I__3399 (
            .O(N__23941),
            .I(N__23872));
    InMux I__3398 (
            .O(N__23940),
            .I(N__23872));
    LocalMux I__3397 (
            .O(N__23931),
            .I(N__23867));
    LocalMux I__3396 (
            .O(N__23922),
            .I(N__23867));
    LocalMux I__3395 (
            .O(N__23913),
            .I(N__23858));
    LocalMux I__3394 (
            .O(N__23904),
            .I(N__23858));
    LocalMux I__3393 (
            .O(N__23895),
            .I(N__23858));
    LocalMux I__3392 (
            .O(N__23886),
            .I(N__23858));
    LocalMux I__3391 (
            .O(N__23881),
            .I(\current_shift_inst.timer_phase.running_i ));
    LocalMux I__3390 (
            .O(N__23872),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv4 I__3389 (
            .O(N__23867),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv12 I__3388 (
            .O(N__23858),
            .I(\current_shift_inst.timer_phase.running_i ));
    InMux I__3387 (
            .O(N__23849),
            .I(N__23846));
    LocalMux I__3386 (
            .O(N__23846),
            .I(N__23843));
    Span4Mux_h I__3385 (
            .O(N__23843),
            .I(N__23840));
    Odrv4 I__3384 (
            .O(N__23840),
            .I(il_max_comp1_c));
    CascadeMux I__3383 (
            .O(N__23837),
            .I(N__23833));
    CascadeMux I__3382 (
            .O(N__23836),
            .I(N__23830));
    InMux I__3381 (
            .O(N__23833),
            .I(N__23827));
    InMux I__3380 (
            .O(N__23830),
            .I(N__23823));
    LocalMux I__3379 (
            .O(N__23827),
            .I(N__23820));
    InMux I__3378 (
            .O(N__23826),
            .I(N__23817));
    LocalMux I__3377 (
            .O(N__23823),
            .I(N__23812));
    Span4Mux_h I__3376 (
            .O(N__23820),
            .I(N__23812));
    LocalMux I__3375 (
            .O(N__23817),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    Odrv4 I__3374 (
            .O(N__23812),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    InMux I__3373 (
            .O(N__23807),
            .I(\current_shift_inst.timer_phase.counter_cry_16 ));
    CascadeMux I__3372 (
            .O(N__23804),
            .I(N__23801));
    InMux I__3371 (
            .O(N__23801),
            .I(N__23796));
    InMux I__3370 (
            .O(N__23800),
            .I(N__23793));
    InMux I__3369 (
            .O(N__23799),
            .I(N__23790));
    LocalMux I__3368 (
            .O(N__23796),
            .I(N__23787));
    LocalMux I__3367 (
            .O(N__23793),
            .I(N__23784));
    LocalMux I__3366 (
            .O(N__23790),
            .I(N__23779));
    Span4Mux_v I__3365 (
            .O(N__23787),
            .I(N__23779));
    Odrv4 I__3364 (
            .O(N__23784),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    Odrv4 I__3363 (
            .O(N__23779),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    InMux I__3362 (
            .O(N__23774),
            .I(\current_shift_inst.timer_phase.counter_cry_17 ));
    InMux I__3361 (
            .O(N__23771),
            .I(N__23764));
    InMux I__3360 (
            .O(N__23770),
            .I(N__23764));
    InMux I__3359 (
            .O(N__23769),
            .I(N__23761));
    LocalMux I__3358 (
            .O(N__23764),
            .I(N__23758));
    LocalMux I__3357 (
            .O(N__23761),
            .I(N__23753));
    Span4Mux_v I__3356 (
            .O(N__23758),
            .I(N__23753));
    Odrv4 I__3355 (
            .O(N__23753),
            .I(\current_shift_inst.timer_phase.counterZ0Z_19 ));
    InMux I__3354 (
            .O(N__23750),
            .I(\current_shift_inst.timer_phase.counter_cry_18 ));
    CascadeMux I__3353 (
            .O(N__23747),
            .I(N__23743));
    CascadeMux I__3352 (
            .O(N__23746),
            .I(N__23740));
    InMux I__3351 (
            .O(N__23743),
            .I(N__23735));
    InMux I__3350 (
            .O(N__23740),
            .I(N__23735));
    LocalMux I__3349 (
            .O(N__23735),
            .I(N__23731));
    InMux I__3348 (
            .O(N__23734),
            .I(N__23728));
    Span4Mux_h I__3347 (
            .O(N__23731),
            .I(N__23725));
    LocalMux I__3346 (
            .O(N__23728),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    Odrv4 I__3345 (
            .O(N__23725),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    InMux I__3344 (
            .O(N__23720),
            .I(\current_shift_inst.timer_phase.counter_cry_19 ));
    CascadeMux I__3343 (
            .O(N__23717),
            .I(N__23713));
    CascadeMux I__3342 (
            .O(N__23716),
            .I(N__23710));
    InMux I__3341 (
            .O(N__23713),
            .I(N__23705));
    InMux I__3340 (
            .O(N__23710),
            .I(N__23705));
    LocalMux I__3339 (
            .O(N__23705),
            .I(N__23701));
    InMux I__3338 (
            .O(N__23704),
            .I(N__23698));
    Span4Mux_h I__3337 (
            .O(N__23701),
            .I(N__23695));
    LocalMux I__3336 (
            .O(N__23698),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    Odrv4 I__3335 (
            .O(N__23695),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    InMux I__3334 (
            .O(N__23690),
            .I(\current_shift_inst.timer_phase.counter_cry_20 ));
    InMux I__3333 (
            .O(N__23687),
            .I(N__23681));
    InMux I__3332 (
            .O(N__23686),
            .I(N__23681));
    LocalMux I__3331 (
            .O(N__23681),
            .I(N__23677));
    InMux I__3330 (
            .O(N__23680),
            .I(N__23674));
    Span4Mux_h I__3329 (
            .O(N__23677),
            .I(N__23671));
    LocalMux I__3328 (
            .O(N__23674),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    Odrv4 I__3327 (
            .O(N__23671),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    InMux I__3326 (
            .O(N__23666),
            .I(\current_shift_inst.timer_phase.counter_cry_21 ));
    InMux I__3325 (
            .O(N__23663),
            .I(N__23656));
    InMux I__3324 (
            .O(N__23662),
            .I(N__23656));
    InMux I__3323 (
            .O(N__23661),
            .I(N__23653));
    LocalMux I__3322 (
            .O(N__23656),
            .I(N__23650));
    LocalMux I__3321 (
            .O(N__23653),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    Odrv4 I__3320 (
            .O(N__23650),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    InMux I__3319 (
            .O(N__23645),
            .I(\current_shift_inst.timer_phase.counter_cry_22 ));
    CascadeMux I__3318 (
            .O(N__23642),
            .I(N__23639));
    InMux I__3317 (
            .O(N__23639),
            .I(N__23635));
    InMux I__3316 (
            .O(N__23638),
            .I(N__23631));
    LocalMux I__3315 (
            .O(N__23635),
            .I(N__23628));
    InMux I__3314 (
            .O(N__23634),
            .I(N__23625));
    LocalMux I__3313 (
            .O(N__23631),
            .I(N__23620));
    Span4Mux_h I__3312 (
            .O(N__23628),
            .I(N__23620));
    LocalMux I__3311 (
            .O(N__23625),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    Odrv4 I__3310 (
            .O(N__23620),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    InMux I__3309 (
            .O(N__23615),
            .I(bfn_8_24_0_));
    CascadeMux I__3308 (
            .O(N__23612),
            .I(N__23608));
    CascadeMux I__3307 (
            .O(N__23611),
            .I(N__23605));
    InMux I__3306 (
            .O(N__23608),
            .I(N__23602));
    InMux I__3305 (
            .O(N__23605),
            .I(N__23598));
    LocalMux I__3304 (
            .O(N__23602),
            .I(N__23595));
    InMux I__3303 (
            .O(N__23601),
            .I(N__23592));
    LocalMux I__3302 (
            .O(N__23598),
            .I(N__23589));
    Span4Mux_h I__3301 (
            .O(N__23595),
            .I(N__23586));
    LocalMux I__3300 (
            .O(N__23592),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    Odrv4 I__3299 (
            .O(N__23589),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    Odrv4 I__3298 (
            .O(N__23586),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    InMux I__3297 (
            .O(N__23579),
            .I(bfn_8_22_0_));
    CascadeMux I__3296 (
            .O(N__23576),
            .I(N__23572));
    InMux I__3295 (
            .O(N__23575),
            .I(N__23568));
    InMux I__3294 (
            .O(N__23572),
            .I(N__23565));
    InMux I__3293 (
            .O(N__23571),
            .I(N__23562));
    LocalMux I__3292 (
            .O(N__23568),
            .I(N__23557));
    LocalMux I__3291 (
            .O(N__23565),
            .I(N__23557));
    LocalMux I__3290 (
            .O(N__23562),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    Odrv4 I__3289 (
            .O(N__23557),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    InMux I__3288 (
            .O(N__23552),
            .I(\current_shift_inst.timer_phase.counter_cry_8 ));
    InMux I__3287 (
            .O(N__23549),
            .I(N__23542));
    InMux I__3286 (
            .O(N__23548),
            .I(N__23542));
    InMux I__3285 (
            .O(N__23547),
            .I(N__23539));
    LocalMux I__3284 (
            .O(N__23542),
            .I(N__23536));
    LocalMux I__3283 (
            .O(N__23539),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    Odrv4 I__3282 (
            .O(N__23536),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    InMux I__3281 (
            .O(N__23531),
            .I(\current_shift_inst.timer_phase.counter_cry_9 ));
    CascadeMux I__3280 (
            .O(N__23528),
            .I(N__23524));
    CascadeMux I__3279 (
            .O(N__23527),
            .I(N__23521));
    InMux I__3278 (
            .O(N__23524),
            .I(N__23515));
    InMux I__3277 (
            .O(N__23521),
            .I(N__23515));
    InMux I__3276 (
            .O(N__23520),
            .I(N__23512));
    LocalMux I__3275 (
            .O(N__23515),
            .I(N__23509));
    LocalMux I__3274 (
            .O(N__23512),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    Odrv4 I__3273 (
            .O(N__23509),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    InMux I__3272 (
            .O(N__23504),
            .I(\current_shift_inst.timer_phase.counter_cry_10 ));
    CascadeMux I__3271 (
            .O(N__23501),
            .I(N__23497));
    CascadeMux I__3270 (
            .O(N__23500),
            .I(N__23494));
    InMux I__3269 (
            .O(N__23497),
            .I(N__23489));
    InMux I__3268 (
            .O(N__23494),
            .I(N__23489));
    LocalMux I__3267 (
            .O(N__23489),
            .I(N__23485));
    InMux I__3266 (
            .O(N__23488),
            .I(N__23482));
    Span4Mux_h I__3265 (
            .O(N__23485),
            .I(N__23479));
    LocalMux I__3264 (
            .O(N__23482),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    Odrv4 I__3263 (
            .O(N__23479),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    InMux I__3262 (
            .O(N__23474),
            .I(\current_shift_inst.timer_phase.counter_cry_11 ));
    CascadeMux I__3261 (
            .O(N__23471),
            .I(N__23468));
    InMux I__3260 (
            .O(N__23468),
            .I(N__23464));
    InMux I__3259 (
            .O(N__23467),
            .I(N__23461));
    LocalMux I__3258 (
            .O(N__23464),
            .I(N__23455));
    LocalMux I__3257 (
            .O(N__23461),
            .I(N__23455));
    InMux I__3256 (
            .O(N__23460),
            .I(N__23452));
    Span4Mux_h I__3255 (
            .O(N__23455),
            .I(N__23449));
    LocalMux I__3254 (
            .O(N__23452),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    Odrv4 I__3253 (
            .O(N__23449),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    InMux I__3252 (
            .O(N__23444),
            .I(\current_shift_inst.timer_phase.counter_cry_12 ));
    InMux I__3251 (
            .O(N__23441),
            .I(N__23435));
    InMux I__3250 (
            .O(N__23440),
            .I(N__23435));
    LocalMux I__3249 (
            .O(N__23435),
            .I(N__23431));
    InMux I__3248 (
            .O(N__23434),
            .I(N__23428));
    Span4Mux_h I__3247 (
            .O(N__23431),
            .I(N__23425));
    LocalMux I__3246 (
            .O(N__23428),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    Odrv4 I__3245 (
            .O(N__23425),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    InMux I__3244 (
            .O(N__23420),
            .I(\current_shift_inst.timer_phase.counter_cry_13 ));
    InMux I__3243 (
            .O(N__23417),
            .I(N__23410));
    InMux I__3242 (
            .O(N__23416),
            .I(N__23410));
    InMux I__3241 (
            .O(N__23415),
            .I(N__23407));
    LocalMux I__3240 (
            .O(N__23410),
            .I(N__23404));
    LocalMux I__3239 (
            .O(N__23407),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    Odrv4 I__3238 (
            .O(N__23404),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    InMux I__3237 (
            .O(N__23399),
            .I(\current_shift_inst.timer_phase.counter_cry_14 ));
    CascadeMux I__3236 (
            .O(N__23396),
            .I(N__23393));
    InMux I__3235 (
            .O(N__23393),
            .I(N__23389));
    InMux I__3234 (
            .O(N__23392),
            .I(N__23385));
    LocalMux I__3233 (
            .O(N__23389),
            .I(N__23382));
    InMux I__3232 (
            .O(N__23388),
            .I(N__23379));
    LocalMux I__3231 (
            .O(N__23385),
            .I(N__23374));
    Span4Mux_h I__3230 (
            .O(N__23382),
            .I(N__23374));
    LocalMux I__3229 (
            .O(N__23379),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    Odrv4 I__3228 (
            .O(N__23374),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    InMux I__3227 (
            .O(N__23369),
            .I(bfn_8_23_0_));
    InMux I__3226 (
            .O(N__23366),
            .I(N__23363));
    LocalMux I__3225 (
            .O(N__23363),
            .I(N__23359));
    InMux I__3224 (
            .O(N__23362),
            .I(N__23356));
    Span4Mux_v I__3223 (
            .O(N__23359),
            .I(N__23350));
    LocalMux I__3222 (
            .O(N__23356),
            .I(N__23350));
    InMux I__3221 (
            .O(N__23355),
            .I(N__23347));
    Odrv4 I__3220 (
            .O(N__23350),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    LocalMux I__3219 (
            .O(N__23347),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    InMux I__3218 (
            .O(N__23342),
            .I(bfn_8_21_0_));
    InMux I__3217 (
            .O(N__23339),
            .I(N__23336));
    LocalMux I__3216 (
            .O(N__23336),
            .I(N__23332));
    InMux I__3215 (
            .O(N__23335),
            .I(N__23329));
    Span4Mux_h I__3214 (
            .O(N__23332),
            .I(N__23323));
    LocalMux I__3213 (
            .O(N__23329),
            .I(N__23323));
    InMux I__3212 (
            .O(N__23328),
            .I(N__23320));
    Odrv4 I__3211 (
            .O(N__23323),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    LocalMux I__3210 (
            .O(N__23320),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    InMux I__3209 (
            .O(N__23315),
            .I(\current_shift_inst.timer_phase.counter_cry_0 ));
    CascadeMux I__3208 (
            .O(N__23312),
            .I(N__23308));
    InMux I__3207 (
            .O(N__23311),
            .I(N__23304));
    InMux I__3206 (
            .O(N__23308),
            .I(N__23301));
    InMux I__3205 (
            .O(N__23307),
            .I(N__23298));
    LocalMux I__3204 (
            .O(N__23304),
            .I(N__23293));
    LocalMux I__3203 (
            .O(N__23301),
            .I(N__23293));
    LocalMux I__3202 (
            .O(N__23298),
            .I(N__23288));
    Span4Mux_v I__3201 (
            .O(N__23293),
            .I(N__23288));
    Odrv4 I__3200 (
            .O(N__23288),
            .I(\current_shift_inst.timer_phase.counterZ0Z_2 ));
    InMux I__3199 (
            .O(N__23285),
            .I(\current_shift_inst.timer_phase.counter_cry_1 ));
    CascadeMux I__3198 (
            .O(N__23282),
            .I(N__23278));
    CascadeMux I__3197 (
            .O(N__23281),
            .I(N__23275));
    InMux I__3196 (
            .O(N__23278),
            .I(N__23269));
    InMux I__3195 (
            .O(N__23275),
            .I(N__23269));
    InMux I__3194 (
            .O(N__23274),
            .I(N__23266));
    LocalMux I__3193 (
            .O(N__23269),
            .I(N__23263));
    LocalMux I__3192 (
            .O(N__23266),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    Odrv4 I__3191 (
            .O(N__23263),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    InMux I__3190 (
            .O(N__23258),
            .I(\current_shift_inst.timer_phase.counter_cry_2 ));
    CascadeMux I__3189 (
            .O(N__23255),
            .I(N__23251));
    CascadeMux I__3188 (
            .O(N__23254),
            .I(N__23248));
    InMux I__3187 (
            .O(N__23251),
            .I(N__23243));
    InMux I__3186 (
            .O(N__23248),
            .I(N__23243));
    LocalMux I__3185 (
            .O(N__23243),
            .I(N__23239));
    InMux I__3184 (
            .O(N__23242),
            .I(N__23236));
    Span4Mux_h I__3183 (
            .O(N__23239),
            .I(N__23233));
    LocalMux I__3182 (
            .O(N__23236),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    Odrv4 I__3181 (
            .O(N__23233),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    InMux I__3180 (
            .O(N__23228),
            .I(\current_shift_inst.timer_phase.counter_cry_3 ));
    InMux I__3179 (
            .O(N__23225),
            .I(N__23219));
    InMux I__3178 (
            .O(N__23224),
            .I(N__23219));
    LocalMux I__3177 (
            .O(N__23219),
            .I(N__23215));
    InMux I__3176 (
            .O(N__23218),
            .I(N__23212));
    Span4Mux_h I__3175 (
            .O(N__23215),
            .I(N__23209));
    LocalMux I__3174 (
            .O(N__23212),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    Odrv4 I__3173 (
            .O(N__23209),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    InMux I__3172 (
            .O(N__23204),
            .I(\current_shift_inst.timer_phase.counter_cry_4 ));
    InMux I__3171 (
            .O(N__23201),
            .I(N__23195));
    InMux I__3170 (
            .O(N__23200),
            .I(N__23195));
    LocalMux I__3169 (
            .O(N__23195),
            .I(N__23191));
    InMux I__3168 (
            .O(N__23194),
            .I(N__23188));
    Span4Mux_h I__3167 (
            .O(N__23191),
            .I(N__23185));
    LocalMux I__3166 (
            .O(N__23188),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    Odrv4 I__3165 (
            .O(N__23185),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    InMux I__3164 (
            .O(N__23180),
            .I(\current_shift_inst.timer_phase.counter_cry_5 ));
    CascadeMux I__3163 (
            .O(N__23177),
            .I(N__23173));
    InMux I__3162 (
            .O(N__23176),
            .I(N__23170));
    InMux I__3161 (
            .O(N__23173),
            .I(N__23167));
    LocalMux I__3160 (
            .O(N__23170),
            .I(N__23162));
    LocalMux I__3159 (
            .O(N__23167),
            .I(N__23162));
    Span4Mux_h I__3158 (
            .O(N__23162),
            .I(N__23158));
    InMux I__3157 (
            .O(N__23161),
            .I(N__23155));
    Span4Mux_h I__3156 (
            .O(N__23158),
            .I(N__23152));
    LocalMux I__3155 (
            .O(N__23155),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    Odrv4 I__3154 (
            .O(N__23152),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    InMux I__3153 (
            .O(N__23147),
            .I(\current_shift_inst.timer_phase.counter_cry_6 ));
    InMux I__3152 (
            .O(N__23144),
            .I(\current_shift_inst.z_5_cry_22 ));
    InMux I__3151 (
            .O(N__23141),
            .I(\current_shift_inst.z_5_cry_23 ));
    InMux I__3150 (
            .O(N__23138),
            .I(bfn_8_20_0_));
    InMux I__3149 (
            .O(N__23135),
            .I(\current_shift_inst.z_5_cry_25 ));
    InMux I__3148 (
            .O(N__23132),
            .I(\current_shift_inst.z_5_cry_26 ));
    InMux I__3147 (
            .O(N__23129),
            .I(\current_shift_inst.z_5_cry_27 ));
    CascadeMux I__3146 (
            .O(N__23126),
            .I(N__23123));
    InMux I__3145 (
            .O(N__23123),
            .I(N__23116));
    InMux I__3144 (
            .O(N__23122),
            .I(N__23116));
    InMux I__3143 (
            .O(N__23121),
            .I(N__23113));
    LocalMux I__3142 (
            .O(N__23116),
            .I(N__23110));
    LocalMux I__3141 (
            .O(N__23113),
            .I(N__23107));
    Odrv12 I__3140 (
            .O(N__23110),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    Odrv4 I__3139 (
            .O(N__23107),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    InMux I__3138 (
            .O(N__23102),
            .I(\current_shift_inst.z_5_cry_28 ));
    InMux I__3137 (
            .O(N__23099),
            .I(N__23096));
    LocalMux I__3136 (
            .O(N__23096),
            .I(N__23081));
    InMux I__3135 (
            .O(N__23095),
            .I(N__23074));
    InMux I__3134 (
            .O(N__23094),
            .I(N__23074));
    InMux I__3133 (
            .O(N__23093),
            .I(N__23074));
    InMux I__3132 (
            .O(N__23092),
            .I(N__23065));
    InMux I__3131 (
            .O(N__23091),
            .I(N__23065));
    InMux I__3130 (
            .O(N__23090),
            .I(N__23065));
    InMux I__3129 (
            .O(N__23089),
            .I(N__23065));
    CascadeMux I__3128 (
            .O(N__23088),
            .I(N__23052));
    CascadeMux I__3127 (
            .O(N__23087),
            .I(N__23047));
    CascadeMux I__3126 (
            .O(N__23086),
            .I(N__23044));
    CascadeMux I__3125 (
            .O(N__23085),
            .I(N__23040));
    CascadeMux I__3124 (
            .O(N__23084),
            .I(N__23037));
    Span4Mux_v I__3123 (
            .O(N__23081),
            .I(N__23020));
    LocalMux I__3122 (
            .O(N__23074),
            .I(N__23020));
    LocalMux I__3121 (
            .O(N__23065),
            .I(N__23020));
    InMux I__3120 (
            .O(N__23064),
            .I(N__23017));
    InMux I__3119 (
            .O(N__23063),
            .I(N__23010));
    InMux I__3118 (
            .O(N__23062),
            .I(N__23010));
    InMux I__3117 (
            .O(N__23061),
            .I(N__23010));
    InMux I__3116 (
            .O(N__23060),
            .I(N__23001));
    InMux I__3115 (
            .O(N__23059),
            .I(N__23001));
    InMux I__3114 (
            .O(N__23058),
            .I(N__23001));
    InMux I__3113 (
            .O(N__23057),
            .I(N__23001));
    CascadeMux I__3112 (
            .O(N__23056),
            .I(N__22998));
    CascadeMux I__3111 (
            .O(N__23055),
            .I(N__22995));
    InMux I__3110 (
            .O(N__23052),
            .I(N__22982));
    InMux I__3109 (
            .O(N__23051),
            .I(N__22982));
    InMux I__3108 (
            .O(N__23050),
            .I(N__22982));
    InMux I__3107 (
            .O(N__23047),
            .I(N__22982));
    InMux I__3106 (
            .O(N__23044),
            .I(N__22982));
    InMux I__3105 (
            .O(N__23043),
            .I(N__22975));
    InMux I__3104 (
            .O(N__23040),
            .I(N__22975));
    InMux I__3103 (
            .O(N__23037),
            .I(N__22975));
    CascadeMux I__3102 (
            .O(N__23036),
            .I(N__22971));
    CascadeMux I__3101 (
            .O(N__23035),
            .I(N__22968));
    CascadeMux I__3100 (
            .O(N__23034),
            .I(N__22964));
    CascadeMux I__3099 (
            .O(N__23033),
            .I(N__22961));
    CascadeMux I__3098 (
            .O(N__23032),
            .I(N__22958));
    CascadeMux I__3097 (
            .O(N__23031),
            .I(N__22954));
    CascadeMux I__3096 (
            .O(N__23030),
            .I(N__22951));
    CascadeMux I__3095 (
            .O(N__23029),
            .I(N__22946));
    CascadeMux I__3094 (
            .O(N__23028),
            .I(N__22943));
    CascadeMux I__3093 (
            .O(N__23027),
            .I(N__22940));
    Span4Mux_s1_h I__3092 (
            .O(N__23020),
            .I(N__22937));
    LocalMux I__3091 (
            .O(N__23017),
            .I(N__22932));
    LocalMux I__3090 (
            .O(N__23010),
            .I(N__22932));
    LocalMux I__3089 (
            .O(N__23001),
            .I(N__22929));
    InMux I__3088 (
            .O(N__22998),
            .I(N__22926));
    InMux I__3087 (
            .O(N__22995),
            .I(N__22921));
    InMux I__3086 (
            .O(N__22994),
            .I(N__22921));
    InMux I__3085 (
            .O(N__22993),
            .I(N__22918));
    LocalMux I__3084 (
            .O(N__22982),
            .I(N__22913));
    LocalMux I__3083 (
            .O(N__22975),
            .I(N__22913));
    InMux I__3082 (
            .O(N__22974),
            .I(N__22906));
    InMux I__3081 (
            .O(N__22971),
            .I(N__22906));
    InMux I__3080 (
            .O(N__22968),
            .I(N__22906));
    InMux I__3079 (
            .O(N__22967),
            .I(N__22897));
    InMux I__3078 (
            .O(N__22964),
            .I(N__22897));
    InMux I__3077 (
            .O(N__22961),
            .I(N__22897));
    InMux I__3076 (
            .O(N__22958),
            .I(N__22897));
    InMux I__3075 (
            .O(N__22957),
            .I(N__22890));
    InMux I__3074 (
            .O(N__22954),
            .I(N__22890));
    InMux I__3073 (
            .O(N__22951),
            .I(N__22890));
    InMux I__3072 (
            .O(N__22950),
            .I(N__22879));
    InMux I__3071 (
            .O(N__22949),
            .I(N__22879));
    InMux I__3070 (
            .O(N__22946),
            .I(N__22879));
    InMux I__3069 (
            .O(N__22943),
            .I(N__22879));
    InMux I__3068 (
            .O(N__22940),
            .I(N__22879));
    Span4Mux_v I__3067 (
            .O(N__22937),
            .I(N__22863));
    Span4Mux_v I__3066 (
            .O(N__22932),
            .I(N__22863));
    Span4Mux_v I__3065 (
            .O(N__22929),
            .I(N__22863));
    LocalMux I__3064 (
            .O(N__22926),
            .I(N__22863));
    LocalMux I__3063 (
            .O(N__22921),
            .I(N__22863));
    LocalMux I__3062 (
            .O(N__22918),
            .I(N__22860));
    Span4Mux_v I__3061 (
            .O(N__22913),
            .I(N__22854));
    LocalMux I__3060 (
            .O(N__22906),
            .I(N__22845));
    LocalMux I__3059 (
            .O(N__22897),
            .I(N__22845));
    LocalMux I__3058 (
            .O(N__22890),
            .I(N__22845));
    LocalMux I__3057 (
            .O(N__22879),
            .I(N__22845));
    CascadeMux I__3056 (
            .O(N__22878),
            .I(N__22842));
    CascadeMux I__3055 (
            .O(N__22877),
            .I(N__22839));
    CascadeMux I__3054 (
            .O(N__22876),
            .I(N__22835));
    CascadeMux I__3053 (
            .O(N__22875),
            .I(N__22832));
    CascadeMux I__3052 (
            .O(N__22874),
            .I(N__22829));
    Span4Mux_h I__3051 (
            .O(N__22863),
            .I(N__22826));
    IoSpan4Mux I__3050 (
            .O(N__22860),
            .I(N__22823));
    InMux I__3049 (
            .O(N__22859),
            .I(N__22820));
    InMux I__3048 (
            .O(N__22858),
            .I(N__22817));
    InMux I__3047 (
            .O(N__22857),
            .I(N__22814));
    Span4Mux_h I__3046 (
            .O(N__22854),
            .I(N__22809));
    Span4Mux_v I__3045 (
            .O(N__22845),
            .I(N__22809));
    InMux I__3044 (
            .O(N__22842),
            .I(N__22804));
    InMux I__3043 (
            .O(N__22839),
            .I(N__22804));
    InMux I__3042 (
            .O(N__22838),
            .I(N__22795));
    InMux I__3041 (
            .O(N__22835),
            .I(N__22795));
    InMux I__3040 (
            .O(N__22832),
            .I(N__22795));
    InMux I__3039 (
            .O(N__22829),
            .I(N__22795));
    Span4Mux_v I__3038 (
            .O(N__22826),
            .I(N__22792));
    Span4Mux_s2_v I__3037 (
            .O(N__22823),
            .I(N__22789));
    LocalMux I__3036 (
            .O(N__22820),
            .I(N__22786));
    LocalMux I__3035 (
            .O(N__22817),
            .I(N__22781));
    LocalMux I__3034 (
            .O(N__22814),
            .I(N__22781));
    Sp12to4 I__3033 (
            .O(N__22809),
            .I(N__22774));
    LocalMux I__3032 (
            .O(N__22804),
            .I(N__22774));
    LocalMux I__3031 (
            .O(N__22795),
            .I(N__22774));
    Sp12to4 I__3030 (
            .O(N__22792),
            .I(N__22771));
    Span4Mux_h I__3029 (
            .O(N__22789),
            .I(N__22768));
    Span4Mux_s2_v I__3028 (
            .O(N__22786),
            .I(N__22765));
    Span4Mux_s2_v I__3027 (
            .O(N__22781),
            .I(N__22762));
    Span12Mux_h I__3026 (
            .O(N__22774),
            .I(N__22759));
    Span12Mux_v I__3025 (
            .O(N__22771),
            .I(N__22754));
    Sp12to4 I__3024 (
            .O(N__22768),
            .I(N__22754));
    Span4Mux_h I__3023 (
            .O(N__22765),
            .I(N__22749));
    Span4Mux_h I__3022 (
            .O(N__22762),
            .I(N__22749));
    Odrv12 I__3021 (
            .O(N__22759),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3020 (
            .O(N__22754),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3019 (
            .O(N__22749),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__3018 (
            .O(N__22742),
            .I(N__22737));
    InMux I__3017 (
            .O(N__22741),
            .I(N__22734));
    InMux I__3016 (
            .O(N__22740),
            .I(N__22731));
    InMux I__3015 (
            .O(N__22737),
            .I(N__22728));
    LocalMux I__3014 (
            .O(N__22734),
            .I(N__22723));
    LocalMux I__3013 (
            .O(N__22731),
            .I(N__22723));
    LocalMux I__3012 (
            .O(N__22728),
            .I(N__22720));
    Odrv12 I__3011 (
            .O(N__22723),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    Odrv4 I__3010 (
            .O(N__22720),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    InMux I__3009 (
            .O(N__22715),
            .I(\current_shift_inst.z_5_cry_29 ));
    InMux I__3008 (
            .O(N__22712),
            .I(\current_shift_inst.z_5_cry_30 ));
    InMux I__3007 (
            .O(N__22709),
            .I(\current_shift_inst.z_5_cry_13 ));
    InMux I__3006 (
            .O(N__22706),
            .I(\current_shift_inst.z_5_cry_14 ));
    InMux I__3005 (
            .O(N__22703),
            .I(\current_shift_inst.z_5_cry_15 ));
    InMux I__3004 (
            .O(N__22700),
            .I(bfn_8_19_0_));
    InMux I__3003 (
            .O(N__22697),
            .I(\current_shift_inst.z_5_cry_17 ));
    InMux I__3002 (
            .O(N__22694),
            .I(\current_shift_inst.z_5_cry_18 ));
    InMux I__3001 (
            .O(N__22691),
            .I(\current_shift_inst.z_5_cry_19 ));
    InMux I__3000 (
            .O(N__22688),
            .I(\current_shift_inst.z_5_cry_20 ));
    InMux I__2999 (
            .O(N__22685),
            .I(\current_shift_inst.z_5_cry_21 ));
    InMux I__2998 (
            .O(N__22682),
            .I(\current_shift_inst.z_5_cry_4 ));
    InMux I__2997 (
            .O(N__22679),
            .I(\current_shift_inst.z_5_cry_5 ));
    InMux I__2996 (
            .O(N__22676),
            .I(\current_shift_inst.z_5_cry_6 ));
    InMux I__2995 (
            .O(N__22673),
            .I(\current_shift_inst.z_5_cry_7 ));
    InMux I__2994 (
            .O(N__22670),
            .I(bfn_8_18_0_));
    InMux I__2993 (
            .O(N__22667),
            .I(\current_shift_inst.z_5_cry_9 ));
    InMux I__2992 (
            .O(N__22664),
            .I(\current_shift_inst.z_5_cry_10 ));
    InMux I__2991 (
            .O(N__22661),
            .I(\current_shift_inst.z_5_cry_11 ));
    InMux I__2990 (
            .O(N__22658),
            .I(\current_shift_inst.z_5_cry_12 ));
    InMux I__2989 (
            .O(N__22655),
            .I(\current_shift_inst.control_input_1_cry_20 ));
    InMux I__2988 (
            .O(N__22652),
            .I(\current_shift_inst.control_input_1_cry_21 ));
    InMux I__2987 (
            .O(N__22649),
            .I(\current_shift_inst.control_input_1_cry_22 ));
    InMux I__2986 (
            .O(N__22646),
            .I(bfn_8_16_0_));
    InMux I__2985 (
            .O(N__22643),
            .I(\current_shift_inst.control_input_1_cry_24 ));
    CascadeMux I__2984 (
            .O(N__22640),
            .I(N__22636));
    InMux I__2983 (
            .O(N__22639),
            .I(N__22631));
    InMux I__2982 (
            .O(N__22636),
            .I(N__22626));
    InMux I__2981 (
            .O(N__22635),
            .I(N__22626));
    InMux I__2980 (
            .O(N__22634),
            .I(N__22623));
    LocalMux I__2979 (
            .O(N__22631),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__2978 (
            .O(N__22626),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__2977 (
            .O(N__22623),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    InMux I__2976 (
            .O(N__22616),
            .I(\current_shift_inst.z_5_cry_1 ));
    InMux I__2975 (
            .O(N__22613),
            .I(N__22608));
    InMux I__2974 (
            .O(N__22612),
            .I(N__22603));
    InMux I__2973 (
            .O(N__22611),
            .I(N__22603));
    LocalMux I__2972 (
            .O(N__22608),
            .I(N__22600));
    LocalMux I__2971 (
            .O(N__22603),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    Odrv4 I__2970 (
            .O(N__22600),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    InMux I__2969 (
            .O(N__22595),
            .I(\current_shift_inst.z_5_cry_2 ));
    InMux I__2968 (
            .O(N__22592),
            .I(\current_shift_inst.z_5_cry_3 ));
    InMux I__2967 (
            .O(N__22589),
            .I(\current_shift_inst.control_input_1_cry_11 ));
    InMux I__2966 (
            .O(N__22586),
            .I(\current_shift_inst.control_input_1_cry_12 ));
    InMux I__2965 (
            .O(N__22583),
            .I(\current_shift_inst.control_input_1_cry_13 ));
    InMux I__2964 (
            .O(N__22580),
            .I(\current_shift_inst.control_input_1_cry_14 ));
    InMux I__2963 (
            .O(N__22577),
            .I(bfn_8_15_0_));
    InMux I__2962 (
            .O(N__22574),
            .I(\current_shift_inst.control_input_1_cry_16 ));
    InMux I__2961 (
            .O(N__22571),
            .I(\current_shift_inst.control_input_1_cry_17 ));
    InMux I__2960 (
            .O(N__22568),
            .I(\current_shift_inst.control_input_1_cry_18 ));
    InMux I__2959 (
            .O(N__22565),
            .I(\current_shift_inst.control_input_1_cry_19 ));
    InMux I__2958 (
            .O(N__22562),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__2957 (
            .O(N__22559),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__2956 (
            .O(N__22556),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__2955 (
            .O(N__22553),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__2954 (
            .O(N__22550),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__2953 (
            .O(N__22547),
            .I(bfn_8_14_0_));
    InMux I__2952 (
            .O(N__22544),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__2951 (
            .O(N__22541),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__2950 (
            .O(N__22538),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__2949 (
            .O(N__22535),
            .I(N__22532));
    LocalMux I__2948 (
            .O(N__22532),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    InMux I__2947 (
            .O(N__22529),
            .I(N__22526));
    LocalMux I__2946 (
            .O(N__22526),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_14 ));
    CascadeMux I__2945 (
            .O(N__22523),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_ ));
    InMux I__2944 (
            .O(N__22520),
            .I(N__22517));
    LocalMux I__2943 (
            .O(N__22517),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    CascadeMux I__2942 (
            .O(N__22514),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__2941 (
            .O(N__22511),
            .I(N__22508));
    LocalMux I__2940 (
            .O(N__22508),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ));
    InMux I__2939 (
            .O(N__22505),
            .I(N__22502));
    LocalMux I__2938 (
            .O(N__22502),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    CascadeMux I__2937 (
            .O(N__22499),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ));
    InMux I__2936 (
            .O(N__22496),
            .I(N__22493));
    LocalMux I__2935 (
            .O(N__22493),
            .I(N__22490));
    Odrv4 I__2934 (
            .O(N__22490),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_5_0 ));
    InMux I__2933 (
            .O(N__22487),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__2932 (
            .O(N__22484),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__2931 (
            .O(N__22481),
            .I(N__22478));
    LocalMux I__2930 (
            .O(N__22478),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    CascadeMux I__2929 (
            .O(N__22475),
            .I(N__22472));
    InMux I__2928 (
            .O(N__22472),
            .I(N__22469));
    LocalMux I__2927 (
            .O(N__22469),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2926 (
            .O(N__22466),
            .I(N__22463));
    InMux I__2925 (
            .O(N__22463),
            .I(N__22460));
    LocalMux I__2924 (
            .O(N__22460),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2923 (
            .O(N__22457),
            .I(N__22454));
    LocalMux I__2922 (
            .O(N__22454),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2921 (
            .O(N__22451),
            .I(N__22448));
    InMux I__2920 (
            .O(N__22448),
            .I(N__22445));
    LocalMux I__2919 (
            .O(N__22445),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2918 (
            .O(N__22442),
            .I(N__22439));
    LocalMux I__2917 (
            .O(N__22439),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2916 (
            .O(N__22436),
            .I(N__22433));
    InMux I__2915 (
            .O(N__22433),
            .I(N__22430));
    LocalMux I__2914 (
            .O(N__22430),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2913 (
            .O(N__22427),
            .I(N__22424));
    LocalMux I__2912 (
            .O(N__22424),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2911 (
            .O(N__22421),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2910 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__2909 (
            .O(N__22415),
            .I(N__22412));
    IoSpan4Mux I__2908 (
            .O(N__22412),
            .I(N__22409));
    Span4Mux_s2_v I__2907 (
            .O(N__22409),
            .I(N__22406));
    Span4Mux_v I__2906 (
            .O(N__22406),
            .I(N__22403));
    Sp12to4 I__2905 (
            .O(N__22403),
            .I(N__22400));
    Span12Mux_h I__2904 (
            .O(N__22400),
            .I(N__22397));
    Odrv12 I__2903 (
            .O(N__22397),
            .I(pwm_output_c));
    InMux I__2902 (
            .O(N__22394),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ));
    InMux I__2901 (
            .O(N__22391),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ));
    CEMux I__2900 (
            .O(N__22388),
            .I(N__22373));
    CEMux I__2899 (
            .O(N__22387),
            .I(N__22373));
    CEMux I__2898 (
            .O(N__22386),
            .I(N__22373));
    CEMux I__2897 (
            .O(N__22385),
            .I(N__22373));
    CEMux I__2896 (
            .O(N__22384),
            .I(N__22373));
    GlobalMux I__2895 (
            .O(N__22373),
            .I(N__22370));
    gio2CtrlBuf I__2894 (
            .O(N__22370),
            .I(\current_shift_inst.timer_phase.N_188_i_g ));
    InMux I__2893 (
            .O(N__22367),
            .I(N__22364));
    LocalMux I__2892 (
            .O(N__22364),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    CascadeMux I__2891 (
            .O(N__22361),
            .I(N__22358));
    InMux I__2890 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__2889 (
            .O(N__22355),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__2888 (
            .O(N__22352),
            .I(N__22349));
    LocalMux I__2887 (
            .O(N__22349),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    CascadeMux I__2886 (
            .O(N__22346),
            .I(N__22343));
    InMux I__2885 (
            .O(N__22343),
            .I(N__22340));
    LocalMux I__2884 (
            .O(N__22340),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2883 (
            .O(N__22337),
            .I(N__22334));
    InMux I__2882 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__2881 (
            .O(N__22331),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__2880 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__2879 (
            .O(N__22325),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2878 (
            .O(N__22322),
            .I(N__22319));
    InMux I__2877 (
            .O(N__22319),
            .I(N__22316));
    LocalMux I__2876 (
            .O(N__22316),
            .I(N__22313));
    Span4Mux_v I__2875 (
            .O(N__22313),
            .I(N__22310));
    Odrv4 I__2874 (
            .O(N__22310),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    InMux I__2873 (
            .O(N__22307),
            .I(N__22304));
    LocalMux I__2872 (
            .O(N__22304),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2871 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__2870 (
            .O(N__22298),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    CascadeMux I__2869 (
            .O(N__22295),
            .I(N__22292));
    InMux I__2868 (
            .O(N__22292),
            .I(N__22289));
    LocalMux I__2867 (
            .O(N__22289),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2866 (
            .O(N__22286),
            .I(N__22283));
    LocalMux I__2865 (
            .O(N__22283),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    CascadeMux I__2864 (
            .O(N__22280),
            .I(N__22277));
    InMux I__2863 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__2862 (
            .O(N__22274),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__2861 (
            .O(N__22271),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ));
    InMux I__2860 (
            .O(N__22268),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ));
    InMux I__2859 (
            .O(N__22265),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ));
    InMux I__2858 (
            .O(N__22262),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ));
    InMux I__2857 (
            .O(N__22259),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ));
    InMux I__2856 (
            .O(N__22256),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ));
    InMux I__2855 (
            .O(N__22253),
            .I(bfn_7_22_0_));
    InMux I__2854 (
            .O(N__22250),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ));
    InMux I__2853 (
            .O(N__22247),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ));
    InMux I__2852 (
            .O(N__22244),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ));
    InMux I__2851 (
            .O(N__22241),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ));
    InMux I__2850 (
            .O(N__22238),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ));
    InMux I__2849 (
            .O(N__22235),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ));
    InMux I__2848 (
            .O(N__22232),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ));
    InMux I__2847 (
            .O(N__22229),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ));
    InMux I__2846 (
            .O(N__22226),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ));
    InMux I__2845 (
            .O(N__22223),
            .I(bfn_7_21_0_));
    InMux I__2844 (
            .O(N__22220),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ));
    InMux I__2843 (
            .O(N__22217),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ));
    InMux I__2842 (
            .O(N__22214),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ));
    InMux I__2841 (
            .O(N__22211),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ));
    InMux I__2840 (
            .O(N__22208),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ));
    InMux I__2839 (
            .O(N__22205),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ));
    InMux I__2838 (
            .O(N__22202),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ));
    InMux I__2837 (
            .O(N__22199),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ));
    InMux I__2836 (
            .O(N__22196),
            .I(bfn_7_20_0_));
    InMux I__2835 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__2834 (
            .O(N__22190),
            .I(N__22187));
    Odrv4 I__2833 (
            .O(N__22187),
            .I(\delay_measurement_inst.delay_hc_reg3lt19_0 ));
    CascadeMux I__2832 (
            .O(N__22184),
            .I(\delay_measurement_inst.delay_hc_reg3lt19_0_cascade_ ));
    CascadeMux I__2831 (
            .O(N__22181),
            .I(N__22178));
    InMux I__2830 (
            .O(N__22178),
            .I(N__22175));
    LocalMux I__2829 (
            .O(N__22175),
            .I(N__22172));
    Span4Mux_v I__2828 (
            .O(N__22172),
            .I(N__22169));
    Odrv4 I__2827 (
            .O(N__22169),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__2826 (
            .O(N__22166),
            .I(N__22163));
    InMux I__2825 (
            .O(N__22163),
            .I(N__22160));
    LocalMux I__2824 (
            .O(N__22160),
            .I(N__22157));
    Span4Mux_v I__2823 (
            .O(N__22157),
            .I(N__22154));
    Odrv4 I__2822 (
            .O(N__22154),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__2821 (
            .O(N__22151),
            .I(N__22144));
    CascadeMux I__2820 (
            .O(N__22150),
            .I(N__22140));
    CascadeMux I__2819 (
            .O(N__22149),
            .I(N__22136));
    InMux I__2818 (
            .O(N__22148),
            .I(N__22121));
    InMux I__2817 (
            .O(N__22147),
            .I(N__22121));
    InMux I__2816 (
            .O(N__22144),
            .I(N__22121));
    InMux I__2815 (
            .O(N__22143),
            .I(N__22121));
    InMux I__2814 (
            .O(N__22140),
            .I(N__22121));
    InMux I__2813 (
            .O(N__22139),
            .I(N__22121));
    InMux I__2812 (
            .O(N__22136),
            .I(N__22121));
    LocalMux I__2811 (
            .O(N__22121),
            .I(N__22118));
    Odrv12 I__2810 (
            .O(N__22118),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    CascadeMux I__2809 (
            .O(N__22115),
            .I(N__22112));
    InMux I__2808 (
            .O(N__22112),
            .I(N__22109));
    LocalMux I__2807 (
            .O(N__22109),
            .I(N__22106));
    Span4Mux_h I__2806 (
            .O(N__22106),
            .I(N__22103));
    Odrv4 I__2805 (
            .O(N__22103),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__2804 (
            .O(N__22100),
            .I(N__22097));
    LocalMux I__2803 (
            .O(N__22097),
            .I(N__22093));
    CascadeMux I__2802 (
            .O(N__22096),
            .I(N__22089));
    Span4Mux_h I__2801 (
            .O(N__22093),
            .I(N__22086));
    CascadeMux I__2800 (
            .O(N__22092),
            .I(N__22082));
    InMux I__2799 (
            .O(N__22089),
            .I(N__22079));
    Span4Mux_v I__2798 (
            .O(N__22086),
            .I(N__22076));
    InMux I__2797 (
            .O(N__22085),
            .I(N__22071));
    InMux I__2796 (
            .O(N__22082),
            .I(N__22071));
    LocalMux I__2795 (
            .O(N__22079),
            .I(clk_10khz_i));
    Odrv4 I__2794 (
            .O(N__22076),
            .I(clk_10khz_i));
    LocalMux I__2793 (
            .O(N__22071),
            .I(clk_10khz_i));
    InMux I__2792 (
            .O(N__22064),
            .I(N__22061));
    LocalMux I__2791 (
            .O(N__22061),
            .I(N__22058));
    Span4Mux_h I__2790 (
            .O(N__22058),
            .I(N__22055));
    Span4Mux_v I__2789 (
            .O(N__22055),
            .I(N__22052));
    Odrv4 I__2788 (
            .O(N__22052),
            .I(clk_10khz_RNIIENAZ0Z2));
    InMux I__2787 (
            .O(N__22049),
            .I(N__22046));
    LocalMux I__2786 (
            .O(N__22046),
            .I(N__22043));
    Odrv4 I__2785 (
            .O(N__22043),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2784 (
            .O(N__22040),
            .I(N__22037));
    LocalMux I__2783 (
            .O(N__22037),
            .I(N__22034));
    Odrv4 I__2782 (
            .O(N__22034),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2781 (
            .O(N__22031),
            .I(N__22028));
    LocalMux I__2780 (
            .O(N__22028),
            .I(N__22025));
    Span4Mux_v I__2779 (
            .O(N__22025),
            .I(N__22022));
    Span4Mux_h I__2778 (
            .O(N__22022),
            .I(N__22019));
    Odrv4 I__2777 (
            .O(N__22019),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2776 (
            .O(N__22016),
            .I(N__22013));
    LocalMux I__2775 (
            .O(N__22013),
            .I(N__22010));
    Span4Mux_v I__2774 (
            .O(N__22010),
            .I(N__22007));
    Span4Mux_h I__2773 (
            .O(N__22007),
            .I(N__22004));
    Odrv4 I__2772 (
            .O(N__22004),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2771 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__2770 (
            .O(N__21998),
            .I(N__21995));
    Span4Mux_v I__2769 (
            .O(N__21995),
            .I(N__21992));
    Odrv4 I__2768 (
            .O(N__21992),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2767 (
            .O(N__21989),
            .I(N__21986));
    InMux I__2766 (
            .O(N__21986),
            .I(N__21983));
    LocalMux I__2765 (
            .O(N__21983),
            .I(N__21980));
    Odrv4 I__2764 (
            .O(N__21980),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__2763 (
            .O(N__21977),
            .I(N__21974));
    InMux I__2762 (
            .O(N__21974),
            .I(N__21971));
    LocalMux I__2761 (
            .O(N__21971),
            .I(N__21968));
    Span4Mux_h I__2760 (
            .O(N__21968),
            .I(N__21965));
    Span4Mux_h I__2759 (
            .O(N__21965),
            .I(N__21962));
    Odrv4 I__2758 (
            .O(N__21962),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2757 (
            .O(N__21959),
            .I(N__21956));
    InMux I__2756 (
            .O(N__21956),
            .I(N__21953));
    LocalMux I__2755 (
            .O(N__21953),
            .I(N__21950));
    Odrv12 I__2754 (
            .O(N__21950),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__2753 (
            .O(N__21947),
            .I(N__21944));
    InMux I__2752 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__2751 (
            .O(N__21941),
            .I(N__21938));
    Span4Mux_v I__2750 (
            .O(N__21938),
            .I(N__21935));
    Odrv4 I__2749 (
            .O(N__21935),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__2748 (
            .O(N__21932),
            .I(N__21928));
    CascadeMux I__2747 (
            .O(N__21931),
            .I(N__21925));
    InMux I__2746 (
            .O(N__21928),
            .I(N__21922));
    InMux I__2745 (
            .O(N__21925),
            .I(N__21919));
    LocalMux I__2744 (
            .O(N__21922),
            .I(N__21916));
    LocalMux I__2743 (
            .O(N__21919),
            .I(N__21913));
    Span4Mux_h I__2742 (
            .O(N__21916),
            .I(N__21910));
    Span4Mux_h I__2741 (
            .O(N__21913),
            .I(N__21907));
    Odrv4 I__2740 (
            .O(N__21910),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    Odrv4 I__2739 (
            .O(N__21907),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2738 (
            .O(N__21902),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2737 (
            .O(N__21899),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    CascadeMux I__2736 (
            .O(N__21896),
            .I(N__21887));
    CascadeMux I__2735 (
            .O(N__21895),
            .I(N__21884));
    CascadeMux I__2734 (
            .O(N__21894),
            .I(N__21881));
    CascadeMux I__2733 (
            .O(N__21893),
            .I(N__21878));
    CascadeMux I__2732 (
            .O(N__21892),
            .I(N__21875));
    CascadeMux I__2731 (
            .O(N__21891),
            .I(N__21872));
    CascadeMux I__2730 (
            .O(N__21890),
            .I(N__21869));
    InMux I__2729 (
            .O(N__21887),
            .I(N__21866));
    InMux I__2728 (
            .O(N__21884),
            .I(N__21863));
    InMux I__2727 (
            .O(N__21881),
            .I(N__21855));
    InMux I__2726 (
            .O(N__21878),
            .I(N__21855));
    InMux I__2725 (
            .O(N__21875),
            .I(N__21850));
    InMux I__2724 (
            .O(N__21872),
            .I(N__21850));
    InMux I__2723 (
            .O(N__21869),
            .I(N__21847));
    LocalMux I__2722 (
            .O(N__21866),
            .I(N__21844));
    LocalMux I__2721 (
            .O(N__21863),
            .I(N__21841));
    InMux I__2720 (
            .O(N__21862),
            .I(N__21836));
    InMux I__2719 (
            .O(N__21861),
            .I(N__21836));
    InMux I__2718 (
            .O(N__21860),
            .I(N__21833));
    LocalMux I__2717 (
            .O(N__21855),
            .I(N__21830));
    LocalMux I__2716 (
            .O(N__21850),
            .I(N__21825));
    LocalMux I__2715 (
            .O(N__21847),
            .I(N__21825));
    Span4Mux_v I__2714 (
            .O(N__21844),
            .I(N__21818));
    Span4Mux_s2_h I__2713 (
            .O(N__21841),
            .I(N__21818));
    LocalMux I__2712 (
            .O(N__21836),
            .I(N__21818));
    LocalMux I__2711 (
            .O(N__21833),
            .I(N__21815));
    Span4Mux_h I__2710 (
            .O(N__21830),
            .I(N__21810));
    Span4Mux_h I__2709 (
            .O(N__21825),
            .I(N__21810));
    Span4Mux_h I__2708 (
            .O(N__21818),
            .I(N__21807));
    Span12Mux_s5_h I__2707 (
            .O(N__21815),
            .I(N__21804));
    Span4Mux_v I__2706 (
            .O(N__21810),
            .I(N__21801));
    Span4Mux_v I__2705 (
            .O(N__21807),
            .I(N__21798));
    Odrv12 I__2704 (
            .O(N__21804),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2703 (
            .O(N__21801),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2702 (
            .O(N__21798),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__2701 (
            .O(N__21791),
            .I(N__21788));
    InMux I__2700 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__2699 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__2698 (
            .O(N__21782),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__2697 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__2696 (
            .O(N__21776),
            .I(N__21773));
    Odrv4 I__2695 (
            .O(N__21773),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2694 (
            .O(N__21770),
            .I(N__21767));
    LocalMux I__2693 (
            .O(N__21767),
            .I(N__21764));
    Span4Mux_v I__2692 (
            .O(N__21764),
            .I(N__21761));
    Span4Mux_h I__2691 (
            .O(N__21761),
            .I(N__21758));
    Odrv4 I__2690 (
            .O(N__21758),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2689 (
            .O(N__21755),
            .I(N__21752));
    LocalMux I__2688 (
            .O(N__21752),
            .I(N__21749));
    Odrv12 I__2687 (
            .O(N__21749),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2686 (
            .O(N__21746),
            .I(N__21743));
    LocalMux I__2685 (
            .O(N__21743),
            .I(N__21740));
    Odrv4 I__2684 (
            .O(N__21740),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2683 (
            .O(N__21737),
            .I(N__21734));
    LocalMux I__2682 (
            .O(N__21734),
            .I(N__21731));
    Span4Mux_h I__2681 (
            .O(N__21731),
            .I(N__21728));
    Odrv4 I__2680 (
            .O(N__21728),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2679 (
            .O(N__21725),
            .I(N__21722));
    LocalMux I__2678 (
            .O(N__21722),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__2677 (
            .O(N__21719),
            .I(N__21715));
    InMux I__2676 (
            .O(N__21718),
            .I(N__21712));
    LocalMux I__2675 (
            .O(N__21715),
            .I(N__21709));
    LocalMux I__2674 (
            .O(N__21712),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    Odrv4 I__2673 (
            .O(N__21709),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2672 (
            .O(N__21704),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2671 (
            .O(N__21701),
            .I(N__21697));
    InMux I__2670 (
            .O(N__21700),
            .I(N__21694));
    LocalMux I__2669 (
            .O(N__21697),
            .I(N__21691));
    LocalMux I__2668 (
            .O(N__21694),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    Odrv4 I__2667 (
            .O(N__21691),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2666 (
            .O(N__21686),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2665 (
            .O(N__21683),
            .I(N__21677));
    InMux I__2664 (
            .O(N__21682),
            .I(N__21677));
    LocalMux I__2663 (
            .O(N__21677),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2662 (
            .O(N__21674),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2661 (
            .O(N__21671),
            .I(N__21668));
    LocalMux I__2660 (
            .O(N__21668),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__2659 (
            .O(N__21665),
            .I(N__21661));
    InMux I__2658 (
            .O(N__21664),
            .I(N__21658));
    LocalMux I__2657 (
            .O(N__21661),
            .I(N__21653));
    LocalMux I__2656 (
            .O(N__21658),
            .I(N__21653));
    Span4Mux_h I__2655 (
            .O(N__21653),
            .I(N__21650));
    Odrv4 I__2654 (
            .O(N__21650),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2653 (
            .O(N__21647),
            .I(bfn_5_12_0_));
    InMux I__2652 (
            .O(N__21644),
            .I(N__21638));
    InMux I__2651 (
            .O(N__21643),
            .I(N__21638));
    LocalMux I__2650 (
            .O(N__21638),
            .I(N__21635));
    Span4Mux_v I__2649 (
            .O(N__21635),
            .I(N__21632));
    Odrv4 I__2648 (
            .O(N__21632),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2647 (
            .O(N__21629),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    CascadeMux I__2646 (
            .O(N__21626),
            .I(N__21622));
    InMux I__2645 (
            .O(N__21625),
            .I(N__21619));
    InMux I__2644 (
            .O(N__21622),
            .I(N__21616));
    LocalMux I__2643 (
            .O(N__21619),
            .I(N__21613));
    LocalMux I__2642 (
            .O(N__21616),
            .I(N__21610));
    Span4Mux_v I__2641 (
            .O(N__21613),
            .I(N__21607));
    Span4Mux_v I__2640 (
            .O(N__21610),
            .I(N__21602));
    Span4Mux_v I__2639 (
            .O(N__21607),
            .I(N__21602));
    Odrv4 I__2638 (
            .O(N__21602),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2637 (
            .O(N__21599),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__2636 (
            .O(N__21596),
            .I(N__21592));
    InMux I__2635 (
            .O(N__21595),
            .I(N__21587));
    InMux I__2634 (
            .O(N__21592),
            .I(N__21587));
    LocalMux I__2633 (
            .O(N__21587),
            .I(N__21584));
    Span4Mux_h I__2632 (
            .O(N__21584),
            .I(N__21581));
    Odrv4 I__2631 (
            .O(N__21581),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2630 (
            .O(N__21578),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2629 (
            .O(N__21575),
            .I(N__21569));
    InMux I__2628 (
            .O(N__21574),
            .I(N__21569));
    LocalMux I__2627 (
            .O(N__21569),
            .I(N__21566));
    Span4Mux_h I__2626 (
            .O(N__21566),
            .I(N__21563));
    Odrv4 I__2625 (
            .O(N__21563),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2624 (
            .O(N__21560),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2623 (
            .O(N__21557),
            .I(N__21551));
    InMux I__2622 (
            .O(N__21556),
            .I(N__21551));
    LocalMux I__2621 (
            .O(N__21551),
            .I(N__21548));
    Span4Mux_h I__2620 (
            .O(N__21548),
            .I(N__21545));
    Odrv4 I__2619 (
            .O(N__21545),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2618 (
            .O(N__21542),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2617 (
            .O(N__21539),
            .I(N__21535));
    InMux I__2616 (
            .O(N__21538),
            .I(N__21532));
    InMux I__2615 (
            .O(N__21535),
            .I(N__21529));
    LocalMux I__2614 (
            .O(N__21532),
            .I(N__21526));
    LocalMux I__2613 (
            .O(N__21529),
            .I(N__21521));
    Span4Mux_v I__2612 (
            .O(N__21526),
            .I(N__21521));
    Odrv4 I__2611 (
            .O(N__21521),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2610 (
            .O(N__21518),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2609 (
            .O(N__21515),
            .I(N__21509));
    InMux I__2608 (
            .O(N__21514),
            .I(N__21509));
    LocalMux I__2607 (
            .O(N__21509),
            .I(N__21506));
    Odrv4 I__2606 (
            .O(N__21506),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2605 (
            .O(N__21503),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2604 (
            .O(N__21500),
            .I(N__21497));
    LocalMux I__2603 (
            .O(N__21497),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    InMux I__2602 (
            .O(N__21494),
            .I(N__21488));
    InMux I__2601 (
            .O(N__21493),
            .I(N__21488));
    LocalMux I__2600 (
            .O(N__21488),
            .I(N__21485));
    Odrv4 I__2599 (
            .O(N__21485),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2598 (
            .O(N__21482),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2597 (
            .O(N__21479),
            .I(N__21476));
    LocalMux I__2596 (
            .O(N__21476),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__2595 (
            .O(N__21473),
            .I(N__21470));
    LocalMux I__2594 (
            .O(N__21470),
            .I(N__21466));
    InMux I__2593 (
            .O(N__21469),
            .I(N__21463));
    Span4Mux_v I__2592 (
            .O(N__21466),
            .I(N__21460));
    LocalMux I__2591 (
            .O(N__21463),
            .I(N__21457));
    Odrv4 I__2590 (
            .O(N__21460),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    Odrv12 I__2589 (
            .O(N__21457),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2588 (
            .O(N__21452),
            .I(bfn_5_11_0_));
    CascadeMux I__2587 (
            .O(N__21449),
            .I(N__21445));
    InMux I__2586 (
            .O(N__21448),
            .I(N__21440));
    InMux I__2585 (
            .O(N__21445),
            .I(N__21440));
    LocalMux I__2584 (
            .O(N__21440),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2583 (
            .O(N__21437),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    CascadeMux I__2582 (
            .O(N__21434),
            .I(N__21431));
    InMux I__2581 (
            .O(N__21431),
            .I(N__21428));
    LocalMux I__2580 (
            .O(N__21428),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__2579 (
            .O(N__21425),
            .I(N__21421));
    InMux I__2578 (
            .O(N__21424),
            .I(N__21418));
    LocalMux I__2577 (
            .O(N__21421),
            .I(N__21415));
    LocalMux I__2576 (
            .O(N__21418),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    Odrv12 I__2575 (
            .O(N__21415),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2574 (
            .O(N__21410),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2573 (
            .O(N__21407),
            .I(N__21401));
    InMux I__2572 (
            .O(N__21406),
            .I(N__21401));
    LocalMux I__2571 (
            .O(N__21401),
            .I(N__21398));
    Odrv4 I__2570 (
            .O(N__21398),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2569 (
            .O(N__21395),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    CascadeMux I__2568 (
            .O(N__21392),
            .I(N__21389));
    InMux I__2567 (
            .O(N__21389),
            .I(N__21386));
    LocalMux I__2566 (
            .O(N__21386),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__2565 (
            .O(N__21383),
            .I(N__21379));
    InMux I__2564 (
            .O(N__21382),
            .I(N__21376));
    LocalMux I__2563 (
            .O(N__21379),
            .I(N__21373));
    LocalMux I__2562 (
            .O(N__21376),
            .I(N__21370));
    Span4Mux_h I__2561 (
            .O(N__21373),
            .I(N__21367));
    Odrv4 I__2560 (
            .O(N__21370),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    Odrv4 I__2559 (
            .O(N__21367),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2558 (
            .O(N__21362),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2557 (
            .O(N__21359),
            .I(N__21356));
    InMux I__2556 (
            .O(N__21356),
            .I(N__21353));
    LocalMux I__2555 (
            .O(N__21353),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__2554 (
            .O(N__21350),
            .I(N__21344));
    InMux I__2553 (
            .O(N__21349),
            .I(N__21344));
    LocalMux I__2552 (
            .O(N__21344),
            .I(N__21340));
    InMux I__2551 (
            .O(N__21343),
            .I(N__21337));
    Span4Mux_s3_h I__2550 (
            .O(N__21340),
            .I(N__21332));
    LocalMux I__2549 (
            .O(N__21337),
            .I(N__21332));
    Span4Mux_v I__2548 (
            .O(N__21332),
            .I(N__21329));
    Odrv4 I__2547 (
            .O(N__21329),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2546 (
            .O(N__21326),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2545 (
            .O(N__21323),
            .I(N__21319));
    InMux I__2544 (
            .O(N__21322),
            .I(N__21316));
    LocalMux I__2543 (
            .O(N__21319),
            .I(N__21310));
    LocalMux I__2542 (
            .O(N__21316),
            .I(N__21310));
    InMux I__2541 (
            .O(N__21315),
            .I(N__21307));
    Span4Mux_v I__2540 (
            .O(N__21310),
            .I(N__21302));
    LocalMux I__2539 (
            .O(N__21307),
            .I(N__21302));
    Span4Mux_h I__2538 (
            .O(N__21302),
            .I(N__21299));
    Odrv4 I__2537 (
            .O(N__21299),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2536 (
            .O(N__21296),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2535 (
            .O(N__21293),
            .I(N__21290));
    LocalMux I__2534 (
            .O(N__21290),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__2533 (
            .O(N__21287),
            .I(N__21283));
    InMux I__2532 (
            .O(N__21286),
            .I(N__21280));
    LocalMux I__2531 (
            .O(N__21283),
            .I(N__21274));
    LocalMux I__2530 (
            .O(N__21280),
            .I(N__21274));
    InMux I__2529 (
            .O(N__21279),
            .I(N__21271));
    Span4Mux_v I__2528 (
            .O(N__21274),
            .I(N__21266));
    LocalMux I__2527 (
            .O(N__21271),
            .I(N__21266));
    Span4Mux_h I__2526 (
            .O(N__21266),
            .I(N__21263));
    Odrv4 I__2525 (
            .O(N__21263),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2524 (
            .O(N__21260),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__2523 (
            .O(N__21257),
            .I(N__21254));
    InMux I__2522 (
            .O(N__21254),
            .I(N__21251));
    LocalMux I__2521 (
            .O(N__21251),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__2520 (
            .O(N__21248),
            .I(N__21244));
    InMux I__2519 (
            .O(N__21247),
            .I(N__21241));
    LocalMux I__2518 (
            .O(N__21244),
            .I(N__21237));
    LocalMux I__2517 (
            .O(N__21241),
            .I(N__21234));
    InMux I__2516 (
            .O(N__21240),
            .I(N__21231));
    Span4Mux_v I__2515 (
            .O(N__21237),
            .I(N__21228));
    Span4Mux_v I__2514 (
            .O(N__21234),
            .I(N__21223));
    LocalMux I__2513 (
            .O(N__21231),
            .I(N__21223));
    Span4Mux_h I__2512 (
            .O(N__21228),
            .I(N__21220));
    Span4Mux_h I__2511 (
            .O(N__21223),
            .I(N__21217));
    Odrv4 I__2510 (
            .O(N__21220),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2509 (
            .O(N__21217),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2508 (
            .O(N__21212),
            .I(bfn_5_10_0_));
    InMux I__2507 (
            .O(N__21209),
            .I(N__21205));
    InMux I__2506 (
            .O(N__21208),
            .I(N__21202));
    LocalMux I__2505 (
            .O(N__21205),
            .I(N__21198));
    LocalMux I__2504 (
            .O(N__21202),
            .I(N__21195));
    InMux I__2503 (
            .O(N__21201),
            .I(N__21192));
    Span4Mux_v I__2502 (
            .O(N__21198),
            .I(N__21189));
    Span4Mux_v I__2501 (
            .O(N__21195),
            .I(N__21184));
    LocalMux I__2500 (
            .O(N__21192),
            .I(N__21184));
    Span4Mux_h I__2499 (
            .O(N__21189),
            .I(N__21181));
    Span4Mux_h I__2498 (
            .O(N__21184),
            .I(N__21178));
    Odrv4 I__2497 (
            .O(N__21181),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2496 (
            .O(N__21178),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2495 (
            .O(N__21173),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    CascadeMux I__2494 (
            .O(N__21170),
            .I(N__21167));
    InMux I__2493 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__2492 (
            .O(N__21164),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2491 (
            .O(N__21161),
            .I(N__21155));
    InMux I__2490 (
            .O(N__21160),
            .I(N__21155));
    LocalMux I__2489 (
            .O(N__21155),
            .I(N__21152));
    Odrv4 I__2488 (
            .O(N__21152),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2487 (
            .O(N__21149),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    CascadeMux I__2486 (
            .O(N__21146),
            .I(N__21143));
    InMux I__2485 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__2484 (
            .O(N__21140),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2483 (
            .O(N__21137),
            .I(N__21133));
    InMux I__2482 (
            .O(N__21136),
            .I(N__21130));
    LocalMux I__2481 (
            .O(N__21133),
            .I(N__21127));
    LocalMux I__2480 (
            .O(N__21130),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    Odrv4 I__2479 (
            .O(N__21127),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2478 (
            .O(N__21122),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__2477 (
            .O(N__21119),
            .I(N__21116));
    InMux I__2476 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__2475 (
            .O(N__21113),
            .I(N__21110));
    Odrv4 I__2474 (
            .O(N__21110),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2473 (
            .O(N__21107),
            .I(N__21101));
    InMux I__2472 (
            .O(N__21106),
            .I(N__21101));
    LocalMux I__2471 (
            .O(N__21101),
            .I(N__21098));
    Odrv4 I__2470 (
            .O(N__21098),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2469 (
            .O(N__21095),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    CascadeMux I__2468 (
            .O(N__21092),
            .I(N__21086));
    InMux I__2467 (
            .O(N__21091),
            .I(N__21077));
    InMux I__2466 (
            .O(N__21090),
            .I(N__21077));
    InMux I__2465 (
            .O(N__21089),
            .I(N__21077));
    InMux I__2464 (
            .O(N__21086),
            .I(N__21074));
    InMux I__2463 (
            .O(N__21085),
            .I(N__21071));
    InMux I__2462 (
            .O(N__21084),
            .I(N__21068));
    LocalMux I__2461 (
            .O(N__21077),
            .I(un2_counter_8));
    LocalMux I__2460 (
            .O(N__21074),
            .I(un2_counter_8));
    LocalMux I__2459 (
            .O(N__21071),
            .I(un2_counter_8));
    LocalMux I__2458 (
            .O(N__21068),
            .I(un2_counter_8));
    InMux I__2457 (
            .O(N__21059),
            .I(N__21051));
    InMux I__2456 (
            .O(N__21058),
            .I(N__21046));
    InMux I__2455 (
            .O(N__21057),
            .I(N__21046));
    InMux I__2454 (
            .O(N__21056),
            .I(N__21043));
    InMux I__2453 (
            .O(N__21055),
            .I(N__21040));
    InMux I__2452 (
            .O(N__21054),
            .I(N__21037));
    LocalMux I__2451 (
            .O(N__21051),
            .I(un2_counter_7));
    LocalMux I__2450 (
            .O(N__21046),
            .I(un2_counter_7));
    LocalMux I__2449 (
            .O(N__21043),
            .I(un2_counter_7));
    LocalMux I__2448 (
            .O(N__21040),
            .I(un2_counter_7));
    LocalMux I__2447 (
            .O(N__21037),
            .I(un2_counter_7));
    InMux I__2446 (
            .O(N__21026),
            .I(N__21018));
    InMux I__2445 (
            .O(N__21025),
            .I(N__21015));
    InMux I__2444 (
            .O(N__21024),
            .I(N__21012));
    InMux I__2443 (
            .O(N__21023),
            .I(N__21005));
    InMux I__2442 (
            .O(N__21022),
            .I(N__21005));
    InMux I__2441 (
            .O(N__21021),
            .I(N__21005));
    LocalMux I__2440 (
            .O(N__21018),
            .I(N__20998));
    LocalMux I__2439 (
            .O(N__21015),
            .I(N__20998));
    LocalMux I__2438 (
            .O(N__21012),
            .I(N__20998));
    LocalMux I__2437 (
            .O(N__21005),
            .I(un2_counter_9));
    Odrv4 I__2436 (
            .O(N__20998),
            .I(un2_counter_9));
    CascadeMux I__2435 (
            .O(N__20993),
            .I(clk_10khz_RNIIENAZ0Z2_cascade_));
    InMux I__2434 (
            .O(N__20990),
            .I(N__20987));
    LocalMux I__2433 (
            .O(N__20987),
            .I(N__20984));
    Span4Mux_v I__2432 (
            .O(N__20984),
            .I(N__20981));
    Odrv4 I__2431 (
            .O(N__20981),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    CascadeMux I__2430 (
            .O(N__20978),
            .I(N__20975));
    InMux I__2429 (
            .O(N__20975),
            .I(N__20972));
    LocalMux I__2428 (
            .O(N__20972),
            .I(N__20969));
    Span4Mux_h I__2427 (
            .O(N__20969),
            .I(N__20966));
    Odrv4 I__2426 (
            .O(N__20966),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__2425 (
            .O(N__20963),
            .I(N__20960));
    InMux I__2424 (
            .O(N__20960),
            .I(N__20957));
    LocalMux I__2423 (
            .O(N__20957),
            .I(N__20954));
    Span4Mux_s2_h I__2422 (
            .O(N__20954),
            .I(N__20951));
    Span4Mux_h I__2421 (
            .O(N__20951),
            .I(N__20948));
    Odrv4 I__2420 (
            .O(N__20948),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2419 (
            .O(N__20945),
            .I(N__20942));
    LocalMux I__2418 (
            .O(N__20942),
            .I(N__20939));
    Span4Mux_h I__2417 (
            .O(N__20939),
            .I(N__20936));
    Odrv4 I__2416 (
            .O(N__20936),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2415 (
            .O(N__20933),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    CascadeMux I__2414 (
            .O(N__20930),
            .I(N__20927));
    InMux I__2413 (
            .O(N__20927),
            .I(N__20924));
    LocalMux I__2412 (
            .O(N__20924),
            .I(N__20921));
    Span4Mux_v I__2411 (
            .O(N__20921),
            .I(N__20918));
    Odrv4 I__2410 (
            .O(N__20918),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2409 (
            .O(N__20915),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    CascadeMux I__2408 (
            .O(N__20912),
            .I(N__20909));
    InMux I__2407 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__2406 (
            .O(N__20906),
            .I(N__20903));
    Span4Mux_v I__2405 (
            .O(N__20903),
            .I(N__20900));
    Odrv4 I__2404 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2403 (
            .O(N__20897),
            .I(N__20893));
    InMux I__2402 (
            .O(N__20896),
            .I(N__20890));
    LocalMux I__2401 (
            .O(N__20893),
            .I(N__20885));
    LocalMux I__2400 (
            .O(N__20890),
            .I(N__20885));
    Span4Mux_h I__2399 (
            .O(N__20885),
            .I(N__20881));
    InMux I__2398 (
            .O(N__20884),
            .I(N__20878));
    Odrv4 I__2397 (
            .O(N__20881),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    LocalMux I__2396 (
            .O(N__20878),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2395 (
            .O(N__20873),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2394 (
            .O(N__20870),
            .I(N__20867));
    LocalMux I__2393 (
            .O(N__20867),
            .I(N__20863));
    InMux I__2392 (
            .O(N__20866),
            .I(N__20860));
    Span4Mux_s3_h I__2391 (
            .O(N__20863),
            .I(N__20854));
    LocalMux I__2390 (
            .O(N__20860),
            .I(N__20854));
    InMux I__2389 (
            .O(N__20859),
            .I(N__20851));
    Span4Mux_h I__2388 (
            .O(N__20854),
            .I(N__20846));
    LocalMux I__2387 (
            .O(N__20851),
            .I(N__20846));
    Span4Mux_v I__2386 (
            .O(N__20846),
            .I(N__20842));
    InMux I__2385 (
            .O(N__20845),
            .I(N__20839));
    Odrv4 I__2384 (
            .O(N__20842),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    LocalMux I__2383 (
            .O(N__20839),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2382 (
            .O(N__20834),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2381 (
            .O(N__20831),
            .I(N__20828));
    LocalMux I__2380 (
            .O(N__20828),
            .I(N__20825));
    Glb2LocalMux I__2379 (
            .O(N__20825),
            .I(N__20822));
    GlobalMux I__2378 (
            .O(N__20822),
            .I(clk_12mhz));
    IoInMux I__2377 (
            .O(N__20819),
            .I(N__20816));
    LocalMux I__2376 (
            .O(N__20816),
            .I(N__20813));
    IoSpan4Mux I__2375 (
            .O(N__20813),
            .I(N__20810));
    Span4Mux_s0_v I__2374 (
            .O(N__20810),
            .I(N__20807));
    Odrv4 I__2373 (
            .O(N__20807),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2372 (
            .O(N__20804),
            .I(N__20800));
    InMux I__2371 (
            .O(N__20803),
            .I(N__20797));
    LocalMux I__2370 (
            .O(N__20800),
            .I(counterZ0Z_4));
    LocalMux I__2369 (
            .O(N__20797),
            .I(counterZ0Z_4));
    InMux I__2368 (
            .O(N__20792),
            .I(N__20788));
    InMux I__2367 (
            .O(N__20791),
            .I(N__20785));
    LocalMux I__2366 (
            .O(N__20788),
            .I(counterZ0Z_3));
    LocalMux I__2365 (
            .O(N__20785),
            .I(counterZ0Z_3));
    InMux I__2364 (
            .O(N__20780),
            .I(N__20776));
    InMux I__2363 (
            .O(N__20779),
            .I(N__20773));
    LocalMux I__2362 (
            .O(N__20776),
            .I(counterZ0Z_5));
    LocalMux I__2361 (
            .O(N__20773),
            .I(counterZ0Z_5));
    InMux I__2360 (
            .O(N__20768),
            .I(N__20764));
    InMux I__2359 (
            .O(N__20767),
            .I(N__20761));
    LocalMux I__2358 (
            .O(N__20764),
            .I(counterZ0Z_6));
    LocalMux I__2357 (
            .O(N__20761),
            .I(counterZ0Z_6));
    CascadeMux I__2356 (
            .O(N__20756),
            .I(un2_counter_5_cascade_));
    CascadeMux I__2355 (
            .O(N__20753),
            .I(N__20750));
    InMux I__2354 (
            .O(N__20750),
            .I(N__20747));
    LocalMux I__2353 (
            .O(N__20747),
            .I(counter_RNO_0Z0Z_12));
    CascadeMux I__2352 (
            .O(N__20744),
            .I(N__20740));
    InMux I__2351 (
            .O(N__20743),
            .I(N__20737));
    InMux I__2350 (
            .O(N__20740),
            .I(N__20734));
    LocalMux I__2349 (
            .O(N__20737),
            .I(counterZ0Z_12));
    LocalMux I__2348 (
            .O(N__20734),
            .I(counterZ0Z_12));
    CascadeMux I__2347 (
            .O(N__20729),
            .I(N__20726));
    InMux I__2346 (
            .O(N__20726),
            .I(N__20723));
    LocalMux I__2345 (
            .O(N__20723),
            .I(counter_RNO_0Z0Z_10));
    CascadeMux I__2344 (
            .O(N__20720),
            .I(N__20716));
    InMux I__2343 (
            .O(N__20719),
            .I(N__20713));
    InMux I__2342 (
            .O(N__20716),
            .I(N__20710));
    LocalMux I__2341 (
            .O(N__20713),
            .I(counterZ0Z_10));
    LocalMux I__2340 (
            .O(N__20710),
            .I(counterZ0Z_10));
    InMux I__2339 (
            .O(N__20705),
            .I(N__20700));
    InMux I__2338 (
            .O(N__20704),
            .I(N__20697));
    InMux I__2337 (
            .O(N__20703),
            .I(N__20694));
    LocalMux I__2336 (
            .O(N__20700),
            .I(counterZ0Z_1));
    LocalMux I__2335 (
            .O(N__20697),
            .I(counterZ0Z_1));
    LocalMux I__2334 (
            .O(N__20694),
            .I(counterZ0Z_1));
    CascadeMux I__2333 (
            .O(N__20687),
            .I(N__20682));
    CascadeMux I__2332 (
            .O(N__20686),
            .I(N__20679));
    InMux I__2331 (
            .O(N__20685),
            .I(N__20673));
    InMux I__2330 (
            .O(N__20682),
            .I(N__20673));
    InMux I__2329 (
            .O(N__20679),
            .I(N__20670));
    InMux I__2328 (
            .O(N__20678),
            .I(N__20667));
    LocalMux I__2327 (
            .O(N__20673),
            .I(counterZ0Z_0));
    LocalMux I__2326 (
            .O(N__20670),
            .I(counterZ0Z_0));
    LocalMux I__2325 (
            .O(N__20667),
            .I(counterZ0Z_0));
    InMux I__2324 (
            .O(N__20660),
            .I(N__20657));
    LocalMux I__2323 (
            .O(N__20657),
            .I(N__20654));
    Odrv12 I__2322 (
            .O(N__20654),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2321 (
            .O(N__20651),
            .I(N__20648));
    LocalMux I__2320 (
            .O(N__20648),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2319 (
            .O(N__20645),
            .I(N__20642));
    LocalMux I__2318 (
            .O(N__20642),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2317 (
            .O(N__20639),
            .I(N__20636));
    LocalMux I__2316 (
            .O(N__20636),
            .I(N__20633));
    Odrv12 I__2315 (
            .O(N__20633),
            .I(counter_RNO_0Z0Z_7));
    InMux I__2314 (
            .O(N__20630),
            .I(N__20627));
    LocalMux I__2313 (
            .O(N__20627),
            .I(N__20623));
    InMux I__2312 (
            .O(N__20626),
            .I(N__20620));
    Odrv4 I__2311 (
            .O(N__20623),
            .I(counterZ0Z_7));
    LocalMux I__2310 (
            .O(N__20620),
            .I(counterZ0Z_7));
    InMux I__2309 (
            .O(N__20615),
            .I(N__20594));
    InMux I__2308 (
            .O(N__20614),
            .I(N__20591));
    InMux I__2307 (
            .O(N__20613),
            .I(N__20574));
    InMux I__2306 (
            .O(N__20612),
            .I(N__20574));
    InMux I__2305 (
            .O(N__20611),
            .I(N__20574));
    InMux I__2304 (
            .O(N__20610),
            .I(N__20574));
    InMux I__2303 (
            .O(N__20609),
            .I(N__20574));
    InMux I__2302 (
            .O(N__20608),
            .I(N__20574));
    InMux I__2301 (
            .O(N__20607),
            .I(N__20574));
    InMux I__2300 (
            .O(N__20606),
            .I(N__20574));
    InMux I__2299 (
            .O(N__20605),
            .I(N__20559));
    InMux I__2298 (
            .O(N__20604),
            .I(N__20559));
    InMux I__2297 (
            .O(N__20603),
            .I(N__20559));
    InMux I__2296 (
            .O(N__20602),
            .I(N__20559));
    InMux I__2295 (
            .O(N__20601),
            .I(N__20559));
    InMux I__2294 (
            .O(N__20600),
            .I(N__20559));
    InMux I__2293 (
            .O(N__20599),
            .I(N__20559));
    InMux I__2292 (
            .O(N__20598),
            .I(N__20548));
    InMux I__2291 (
            .O(N__20597),
            .I(N__20548));
    LocalMux I__2290 (
            .O(N__20594),
            .I(N__20545));
    LocalMux I__2289 (
            .O(N__20591),
            .I(N__20540));
    LocalMux I__2288 (
            .O(N__20574),
            .I(N__20540));
    LocalMux I__2287 (
            .O(N__20559),
            .I(N__20537));
    InMux I__2286 (
            .O(N__20558),
            .I(N__20532));
    InMux I__2285 (
            .O(N__20557),
            .I(N__20532));
    CascadeMux I__2284 (
            .O(N__20556),
            .I(N__20526));
    CascadeMux I__2283 (
            .O(N__20555),
            .I(N__20523));
    CascadeMux I__2282 (
            .O(N__20554),
            .I(N__20520));
    CascadeMux I__2281 (
            .O(N__20553),
            .I(N__20517));
    LocalMux I__2280 (
            .O(N__20548),
            .I(N__20510));
    Span4Mux_v I__2279 (
            .O(N__20545),
            .I(N__20503));
    Span4Mux_v I__2278 (
            .O(N__20540),
            .I(N__20503));
    Span4Mux_v I__2277 (
            .O(N__20537),
            .I(N__20503));
    LocalMux I__2276 (
            .O(N__20532),
            .I(N__20500));
    InMux I__2275 (
            .O(N__20531),
            .I(N__20493));
    InMux I__2274 (
            .O(N__20530),
            .I(N__20493));
    InMux I__2273 (
            .O(N__20529),
            .I(N__20493));
    InMux I__2272 (
            .O(N__20526),
            .I(N__20488));
    InMux I__2271 (
            .O(N__20523),
            .I(N__20488));
    InMux I__2270 (
            .O(N__20520),
            .I(N__20483));
    InMux I__2269 (
            .O(N__20517),
            .I(N__20483));
    InMux I__2268 (
            .O(N__20516),
            .I(N__20474));
    InMux I__2267 (
            .O(N__20515),
            .I(N__20474));
    InMux I__2266 (
            .O(N__20514),
            .I(N__20474));
    InMux I__2265 (
            .O(N__20513),
            .I(N__20474));
    Span4Mux_v I__2264 (
            .O(N__20510),
            .I(N__20471));
    Span4Mux_v I__2263 (
            .O(N__20503),
            .I(N__20466));
    Span4Mux_s1_h I__2262 (
            .O(N__20500),
            .I(N__20466));
    LocalMux I__2261 (
            .O(N__20493),
            .I(N__20463));
    LocalMux I__2260 (
            .O(N__20488),
            .I(N_19_1));
    LocalMux I__2259 (
            .O(N__20483),
            .I(N_19_1));
    LocalMux I__2258 (
            .O(N__20474),
            .I(N_19_1));
    Odrv4 I__2257 (
            .O(N__20471),
            .I(N_19_1));
    Odrv4 I__2256 (
            .O(N__20466),
            .I(N_19_1));
    Odrv12 I__2255 (
            .O(N__20463),
            .I(N_19_1));
    InMux I__2254 (
            .O(N__20450),
            .I(N__20432));
    InMux I__2253 (
            .O(N__20449),
            .I(N__20432));
    InMux I__2252 (
            .O(N__20448),
            .I(N__20432));
    InMux I__2251 (
            .O(N__20447),
            .I(N__20432));
    InMux I__2250 (
            .O(N__20446),
            .I(N__20432));
    InMux I__2249 (
            .O(N__20445),
            .I(N__20432));
    LocalMux I__2248 (
            .O(N__20432),
            .I(N__20427));
    InMux I__2247 (
            .O(N__20431),
            .I(N__20422));
    InMux I__2246 (
            .O(N__20430),
            .I(N__20422));
    Span4Mux_v I__2245 (
            .O(N__20427),
            .I(N__20417));
    LocalMux I__2244 (
            .O(N__20422),
            .I(N__20414));
    InMux I__2243 (
            .O(N__20421),
            .I(N__20409));
    InMux I__2242 (
            .O(N__20420),
            .I(N__20409));
    Odrv4 I__2241 (
            .O(N__20417),
            .I(\pwm_generator_inst.N_17 ));
    Odrv12 I__2240 (
            .O(N__20414),
            .I(\pwm_generator_inst.N_17 ));
    LocalMux I__2239 (
            .O(N__20409),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2238 (
            .O(N__20402),
            .I(N__20392));
    InMux I__2237 (
            .O(N__20401),
            .I(N__20392));
    CascadeMux I__2236 (
            .O(N__20400),
            .I(N__20389));
    CascadeMux I__2235 (
            .O(N__20399),
            .I(N__20386));
    CascadeMux I__2234 (
            .O(N__20398),
            .I(N__20383));
    CascadeMux I__2233 (
            .O(N__20397),
            .I(N__20380));
    LocalMux I__2232 (
            .O(N__20392),
            .I(N__20375));
    InMux I__2231 (
            .O(N__20389),
            .I(N__20362));
    InMux I__2230 (
            .O(N__20386),
            .I(N__20362));
    InMux I__2229 (
            .O(N__20383),
            .I(N__20362));
    InMux I__2228 (
            .O(N__20380),
            .I(N__20362));
    InMux I__2227 (
            .O(N__20379),
            .I(N__20362));
    InMux I__2226 (
            .O(N__20378),
            .I(N__20362));
    Span4Mux_v I__2225 (
            .O(N__20375),
            .I(N__20357));
    LocalMux I__2224 (
            .O(N__20362),
            .I(N__20354));
    InMux I__2223 (
            .O(N__20361),
            .I(N__20349));
    InMux I__2222 (
            .O(N__20360),
            .I(N__20349));
    Odrv4 I__2221 (
            .O(N__20357),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2220 (
            .O(N__20354),
            .I(\pwm_generator_inst.N_16 ));
    LocalMux I__2219 (
            .O(N__20349),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__2218 (
            .O(N__20342),
            .I(N__20339));
    LocalMux I__2217 (
            .O(N__20339),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    CascadeMux I__2216 (
            .O(N__20336),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2215 (
            .O(N__20333),
            .I(N__20330));
    LocalMux I__2214 (
            .O(N__20330),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2213 (
            .O(N__20327),
            .I(N__20324));
    LocalMux I__2212 (
            .O(N__20324),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2211 (
            .O(N__20321),
            .I(un5_counter_cry_9));
    InMux I__2210 (
            .O(N__20318),
            .I(un5_counter_cry_10));
    InMux I__2209 (
            .O(N__20315),
            .I(un5_counter_cry_11));
    InMux I__2208 (
            .O(N__20312),
            .I(N__20308));
    InMux I__2207 (
            .O(N__20311),
            .I(N__20305));
    LocalMux I__2206 (
            .O(N__20308),
            .I(N__20302));
    LocalMux I__2205 (
            .O(N__20305),
            .I(counterZ0Z_11));
    Odrv4 I__2204 (
            .O(N__20302),
            .I(counterZ0Z_11));
    InMux I__2203 (
            .O(N__20297),
            .I(N__20293));
    InMux I__2202 (
            .O(N__20296),
            .I(N__20290));
    LocalMux I__2201 (
            .O(N__20293),
            .I(counterZ0Z_9));
    LocalMux I__2200 (
            .O(N__20290),
            .I(counterZ0Z_9));
    InMux I__2199 (
            .O(N__20285),
            .I(N__20281));
    InMux I__2198 (
            .O(N__20284),
            .I(N__20278));
    LocalMux I__2197 (
            .O(N__20281),
            .I(N__20275));
    LocalMux I__2196 (
            .O(N__20278),
            .I(counterZ0Z_8));
    Odrv4 I__2195 (
            .O(N__20275),
            .I(counterZ0Z_8));
    InMux I__2194 (
            .O(N__20270),
            .I(N__20266));
    InMux I__2193 (
            .O(N__20269),
            .I(N__20263));
    LocalMux I__2192 (
            .O(N__20266),
            .I(N__20260));
    LocalMux I__2191 (
            .O(N__20263),
            .I(counterZ0Z_2));
    Odrv4 I__2190 (
            .O(N__20260),
            .I(counterZ0Z_2));
    InMux I__2189 (
            .O(N__20255),
            .I(N__20252));
    LocalMux I__2188 (
            .O(N__20252),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__2187 (
            .O(N__20249),
            .I(N__20246));
    LocalMux I__2186 (
            .O(N__20246),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2185 (
            .O(N__20243),
            .I(N__20240));
    LocalMux I__2184 (
            .O(N__20240),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__2183 (
            .O(N__20237),
            .I(N__20234));
    LocalMux I__2182 (
            .O(N__20234),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2181 (
            .O(N__20231),
            .I(un5_counter_cry_1));
    InMux I__2180 (
            .O(N__20228),
            .I(un5_counter_cry_2));
    InMux I__2179 (
            .O(N__20225),
            .I(un5_counter_cry_3));
    InMux I__2178 (
            .O(N__20222),
            .I(un5_counter_cry_4));
    InMux I__2177 (
            .O(N__20219),
            .I(un5_counter_cry_5));
    InMux I__2176 (
            .O(N__20216),
            .I(un5_counter_cry_6));
    InMux I__2175 (
            .O(N__20213),
            .I(un5_counter_cry_7));
    InMux I__2174 (
            .O(N__20210),
            .I(bfn_4_6_0_));
    CascadeMux I__2173 (
            .O(N__20207),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ));
    InMux I__2172 (
            .O(N__20204),
            .I(N__20201));
    LocalMux I__2171 (
            .O(N__20201),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2170 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__2169 (
            .O(N__20195),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    CascadeMux I__2168 (
            .O(N__20192),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    InMux I__2167 (
            .O(N__20189),
            .I(N__20186));
    LocalMux I__2166 (
            .O(N__20186),
            .I(N__20183));
    Odrv4 I__2165 (
            .O(N__20183),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    CascadeMux I__2164 (
            .O(N__20180),
            .I(N__20177));
    InMux I__2163 (
            .O(N__20177),
            .I(N__20174));
    LocalMux I__2162 (
            .O(N__20174),
            .I(N__20171));
    Odrv4 I__2161 (
            .O(N__20171),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__2160 (
            .O(N__20168),
            .I(N__20164));
    InMux I__2159 (
            .O(N__20167),
            .I(N__20160));
    LocalMux I__2158 (
            .O(N__20164),
            .I(N__20157));
    InMux I__2157 (
            .O(N__20163),
            .I(N__20154));
    LocalMux I__2156 (
            .O(N__20160),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__2155 (
            .O(N__20157),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2154 (
            .O(N__20154),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__2153 (
            .O(N__20147),
            .I(N__20144));
    LocalMux I__2152 (
            .O(N__20144),
            .I(N__20141));
    Span4Mux_v I__2151 (
            .O(N__20141),
            .I(N__20137));
    InMux I__2150 (
            .O(N__20140),
            .I(N__20134));
    Odrv4 I__2149 (
            .O(N__20137),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    LocalMux I__2148 (
            .O(N__20134),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    CascadeMux I__2147 (
            .O(N__20129),
            .I(N__20126));
    InMux I__2146 (
            .O(N__20126),
            .I(N__20123));
    LocalMux I__2145 (
            .O(N__20123),
            .I(N__20120));
    Span4Mux_h I__2144 (
            .O(N__20120),
            .I(N__20117));
    Span4Mux_v I__2143 (
            .O(N__20117),
            .I(N__20114));
    Odrv4 I__2142 (
            .O(N__20114),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__2141 (
            .O(N__20111),
            .I(N__20108));
    LocalMux I__2140 (
            .O(N__20108),
            .I(N__20105));
    Span4Mux_h I__2139 (
            .O(N__20105),
            .I(N__20102));
    Odrv4 I__2138 (
            .O(N__20102),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__2137 (
            .O(N__20099),
            .I(N__20094));
    InMux I__2136 (
            .O(N__20098),
            .I(N__20091));
    InMux I__2135 (
            .O(N__20097),
            .I(N__20088));
    LocalMux I__2134 (
            .O(N__20094),
            .I(N__20085));
    LocalMux I__2133 (
            .O(N__20091),
            .I(N__20082));
    LocalMux I__2132 (
            .O(N__20088),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__2131 (
            .O(N__20085),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__2130 (
            .O(N__20082),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__2129 (
            .O(N__20075),
            .I(N__20072));
    LocalMux I__2128 (
            .O(N__20072),
            .I(N__20069));
    Span4Mux_h I__2127 (
            .O(N__20069),
            .I(N__20065));
    InMux I__2126 (
            .O(N__20068),
            .I(N__20062));
    Odrv4 I__2125 (
            .O(N__20065),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    LocalMux I__2124 (
            .O(N__20062),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    CascadeMux I__2123 (
            .O(N__20057),
            .I(N__20054));
    InMux I__2122 (
            .O(N__20054),
            .I(N__20051));
    LocalMux I__2121 (
            .O(N__20051),
            .I(N__20048));
    Span4Mux_v I__2120 (
            .O(N__20048),
            .I(N__20045));
    Odrv4 I__2119 (
            .O(N__20045),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    CascadeMux I__2118 (
            .O(N__20042),
            .I(N__20037));
    InMux I__2117 (
            .O(N__20041),
            .I(N__20027));
    InMux I__2116 (
            .O(N__20040),
            .I(N__20024));
    InMux I__2115 (
            .O(N__20037),
            .I(N__20021));
    InMux I__2114 (
            .O(N__20036),
            .I(N__20012));
    InMux I__2113 (
            .O(N__20035),
            .I(N__20012));
    InMux I__2112 (
            .O(N__20034),
            .I(N__20012));
    InMux I__2111 (
            .O(N__20033),
            .I(N__20012));
    InMux I__2110 (
            .O(N__20032),
            .I(N__20007));
    InMux I__2109 (
            .O(N__20031),
            .I(N__20007));
    InMux I__2108 (
            .O(N__20030),
            .I(N__20004));
    LocalMux I__2107 (
            .O(N__20027),
            .I(N__19997));
    LocalMux I__2106 (
            .O(N__20024),
            .I(N__19997));
    LocalMux I__2105 (
            .O(N__20021),
            .I(N__19997));
    LocalMux I__2104 (
            .O(N__20012),
            .I(N__19990));
    LocalMux I__2103 (
            .O(N__20007),
            .I(N__19990));
    LocalMux I__2102 (
            .O(N__20004),
            .I(N__19987));
    Span4Mux_v I__2101 (
            .O(N__19997),
            .I(N__19984));
    InMux I__2100 (
            .O(N__19996),
            .I(N__19979));
    InMux I__2099 (
            .O(N__19995),
            .I(N__19979));
    Span4Mux_v I__2098 (
            .O(N__19990),
            .I(N__19974));
    Span4Mux_v I__2097 (
            .O(N__19987),
            .I(N__19974));
    Odrv4 I__2096 (
            .O(N__19984),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2095 (
            .O(N__19979),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2094 (
            .O(N__19974),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2093 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__2092 (
            .O(N__19964),
            .I(N__19961));
    Odrv12 I__2091 (
            .O(N__19961),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__2090 (
            .O(N__19958),
            .I(N__19955));
    LocalMux I__2089 (
            .O(N__19955),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2088 (
            .O(N__19952),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    CascadeMux I__2087 (
            .O(N__19949),
            .I(N__19946));
    InMux I__2086 (
            .O(N__19946),
            .I(N__19943));
    LocalMux I__2085 (
            .O(N__19943),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    CascadeMux I__2084 (
            .O(N__19940),
            .I(N__19937));
    InMux I__2083 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__2082 (
            .O(N__19934),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2081 (
            .O(N__19931),
            .I(bfn_3_9_0_));
    InMux I__2080 (
            .O(N__19928),
            .I(N__19925));
    LocalMux I__2079 (
            .O(N__19925),
            .I(N__19922));
    Odrv4 I__2078 (
            .O(N__19922),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    CascadeMux I__2077 (
            .O(N__19919),
            .I(N__19916));
    InMux I__2076 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__2075 (
            .O(N__19913),
            .I(N__19910));
    Span4Mux_h I__2074 (
            .O(N__19910),
            .I(N__19907));
    Odrv4 I__2073 (
            .O(N__19907),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2072 (
            .O(N__19904),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    CascadeMux I__2071 (
            .O(N__19901),
            .I(N__19898));
    InMux I__2070 (
            .O(N__19898),
            .I(N__19895));
    LocalMux I__2069 (
            .O(N__19895),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2068 (
            .O(N__19892),
            .I(N__19882));
    InMux I__2067 (
            .O(N__19891),
            .I(N__19877));
    InMux I__2066 (
            .O(N__19890),
            .I(N__19877));
    InMux I__2065 (
            .O(N__19889),
            .I(N__19872));
    InMux I__2064 (
            .O(N__19888),
            .I(N__19872));
    InMux I__2063 (
            .O(N__19887),
            .I(N__19867));
    InMux I__2062 (
            .O(N__19886),
            .I(N__19867));
    InMux I__2061 (
            .O(N__19885),
            .I(N__19864));
    LocalMux I__2060 (
            .O(N__19882),
            .I(N__19858));
    LocalMux I__2059 (
            .O(N__19877),
            .I(N__19858));
    LocalMux I__2058 (
            .O(N__19872),
            .I(N__19855));
    LocalMux I__2057 (
            .O(N__19867),
            .I(N__19850));
    LocalMux I__2056 (
            .O(N__19864),
            .I(N__19850));
    InMux I__2055 (
            .O(N__19863),
            .I(N__19847));
    Span12Mux_s8_v I__2054 (
            .O(N__19858),
            .I(N__19844));
    Span4Mux_v I__2053 (
            .O(N__19855),
            .I(N__19839));
    Span4Mux_s3_h I__2052 (
            .O(N__19850),
            .I(N__19839));
    LocalMux I__2051 (
            .O(N__19847),
            .I(N__19836));
    Odrv12 I__2050 (
            .O(N__19844),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    Odrv4 I__2049 (
            .O(N__19839),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    Odrv12 I__2048 (
            .O(N__19836),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    InMux I__2047 (
            .O(N__19829),
            .I(N__19823));
    InMux I__2046 (
            .O(N__19828),
            .I(N__19816));
    InMux I__2045 (
            .O(N__19827),
            .I(N__19816));
    InMux I__2044 (
            .O(N__19826),
            .I(N__19816));
    LocalMux I__2043 (
            .O(N__19823),
            .I(N__19810));
    LocalMux I__2042 (
            .O(N__19816),
            .I(N__19807));
    InMux I__2041 (
            .O(N__19815),
            .I(N__19802));
    InMux I__2040 (
            .O(N__19814),
            .I(N__19802));
    InMux I__2039 (
            .O(N__19813),
            .I(N__19799));
    Span4Mux_v I__2038 (
            .O(N__19810),
            .I(N__19794));
    Span4Mux_s2_h I__2037 (
            .O(N__19807),
            .I(N__19794));
    LocalMux I__2036 (
            .O(N__19802),
            .I(N__19791));
    LocalMux I__2035 (
            .O(N__19799),
            .I(N__19788));
    Span4Mux_v I__2034 (
            .O(N__19794),
            .I(N__19785));
    Span4Mux_v I__2033 (
            .O(N__19791),
            .I(N__19780));
    Span4Mux_s3_h I__2032 (
            .O(N__19788),
            .I(N__19780));
    Odrv4 I__2031 (
            .O(N__19785),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2030 (
            .O(N__19780),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2029 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__2028 (
            .O(N__19772),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2027 (
            .O(N__19769),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__2026 (
            .O(N__19766),
            .I(N__19763));
    LocalMux I__2025 (
            .O(N__19763),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__2024 (
            .O(N__19760),
            .I(N__19757));
    InMux I__2023 (
            .O(N__19757),
            .I(N__19754));
    LocalMux I__2022 (
            .O(N__19754),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2021 (
            .O(N__19751),
            .I(N__19748));
    LocalMux I__2020 (
            .O(N__19748),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    CascadeMux I__2019 (
            .O(N__19745),
            .I(N__19742));
    InMux I__2018 (
            .O(N__19742),
            .I(N__19739));
    LocalMux I__2017 (
            .O(N__19739),
            .I(N__19736));
    Odrv4 I__2016 (
            .O(N__19736),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2015 (
            .O(N__19733),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__2014 (
            .O(N__19730),
            .I(N__19727));
    LocalMux I__2013 (
            .O(N__19727),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__2012 (
            .O(N__19724),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__2011 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__2010 (
            .O(N__19718),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2009 (
            .O(N__19715),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__2008 (
            .O(N__19712),
            .I(N__19709));
    LocalMux I__2007 (
            .O(N__19709),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__2006 (
            .O(N__19706),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__2005 (
            .O(N__19703),
            .I(N__19700));
    LocalMux I__2004 (
            .O(N__19700),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__2003 (
            .O(N__19697),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__2002 (
            .O(N__19694),
            .I(N__19691));
    LocalMux I__2001 (
            .O(N__19691),
            .I(N__19688));
    Odrv4 I__2000 (
            .O(N__19688),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__1999 (
            .O(N__19685),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__1998 (
            .O(N__19682),
            .I(N__19679));
    LocalMux I__1997 (
            .O(N__19679),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1996 (
            .O(N__19676),
            .I(N__19669));
    CascadeMux I__1995 (
            .O(N__19675),
            .I(N__19666));
    CascadeMux I__1994 (
            .O(N__19674),
            .I(N__19662));
    CascadeMux I__1993 (
            .O(N__19673),
            .I(N__19658));
    InMux I__1992 (
            .O(N__19672),
            .I(N__19654));
    LocalMux I__1991 (
            .O(N__19669),
            .I(N__19651));
    InMux I__1990 (
            .O(N__19666),
            .I(N__19638));
    InMux I__1989 (
            .O(N__19665),
            .I(N__19638));
    InMux I__1988 (
            .O(N__19662),
            .I(N__19638));
    InMux I__1987 (
            .O(N__19661),
            .I(N__19638));
    InMux I__1986 (
            .O(N__19658),
            .I(N__19638));
    InMux I__1985 (
            .O(N__19657),
            .I(N__19638));
    LocalMux I__1984 (
            .O(N__19654),
            .I(N__19631));
    Span4Mux_v I__1983 (
            .O(N__19651),
            .I(N__19631));
    LocalMux I__1982 (
            .O(N__19638),
            .I(N__19631));
    Span4Mux_v I__1981 (
            .O(N__19631),
            .I(N__19628));
    Odrv4 I__1980 (
            .O(N__19628),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1979 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__1978 (
            .O(N__19622),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1977 (
            .O(N__19619),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1976 (
            .O(N__19616),
            .I(N__19613));
    LocalMux I__1975 (
            .O(N__19613),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1974 (
            .O(N__19610),
            .I(N__19607));
    LocalMux I__1973 (
            .O(N__19607),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1972 (
            .O(N__19604),
            .I(bfn_2_13_0_));
    InMux I__1971 (
            .O(N__19601),
            .I(N__19598));
    LocalMux I__1970 (
            .O(N__19598),
            .I(N__19595));
    Span4Mux_s1_v I__1969 (
            .O(N__19595),
            .I(N__19592));
    Odrv4 I__1968 (
            .O(N__19592),
            .I(N_32_i_i));
    InMux I__1967 (
            .O(N__19589),
            .I(N__19586));
    LocalMux I__1966 (
            .O(N__19586),
            .I(N__19583));
    Odrv4 I__1965 (
            .O(N__19583),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__1964 (
            .O(N__19580),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__1963 (
            .O(N__19577),
            .I(N__19572));
    InMux I__1962 (
            .O(N__19576),
            .I(N__19567));
    InMux I__1961 (
            .O(N__19575),
            .I(N__19567));
    LocalMux I__1960 (
            .O(N__19572),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1959 (
            .O(N__19567),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__1958 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__1957 (
            .O(N__19559),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__1956 (
            .O(N__19556),
            .I(N__19552));
    InMux I__1955 (
            .O(N__19555),
            .I(N__19548));
    LocalMux I__1954 (
            .O(N__19552),
            .I(N__19545));
    InMux I__1953 (
            .O(N__19551),
            .I(N__19542));
    LocalMux I__1952 (
            .O(N__19548),
            .I(pwm_duty_input_3));
    Odrv4 I__1951 (
            .O(N__19545),
            .I(pwm_duty_input_3));
    LocalMux I__1950 (
            .O(N__19542),
            .I(pwm_duty_input_3));
    CascadeMux I__1949 (
            .O(N__19535),
            .I(N__19532));
    InMux I__1948 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__1947 (
            .O(N__19529),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__1946 (
            .O(N__19526),
            .I(N__19522));
    InMux I__1945 (
            .O(N__19525),
            .I(N__19519));
    LocalMux I__1944 (
            .O(N__19522),
            .I(N__19515));
    LocalMux I__1943 (
            .O(N__19519),
            .I(N__19512));
    InMux I__1942 (
            .O(N__19518),
            .I(N__19509));
    Span4Mux_v I__1941 (
            .O(N__19515),
            .I(N__19504));
    Span4Mux_v I__1940 (
            .O(N__19512),
            .I(N__19504));
    LocalMux I__1939 (
            .O(N__19509),
            .I(pwm_duty_input_4));
    Odrv4 I__1938 (
            .O(N__19504),
            .I(pwm_duty_input_4));
    InMux I__1937 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__1936 (
            .O(N__19496),
            .I(N__19493));
    Span4Mux_v I__1935 (
            .O(N__19493),
            .I(N__19490));
    Odrv4 I__1934 (
            .O(N__19490),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__1933 (
            .O(N__19487),
            .I(N__19484));
    InMux I__1932 (
            .O(N__19484),
            .I(N__19481));
    LocalMux I__1931 (
            .O(N__19481),
            .I(N__19478));
    Span4Mux_h I__1930 (
            .O(N__19478),
            .I(N__19475));
    Odrv4 I__1929 (
            .O(N__19475),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    InMux I__1928 (
            .O(N__19472),
            .I(N__19469));
    LocalMux I__1927 (
            .O(N__19469),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1926 (
            .O(N__19466),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1925 (
            .O(N__19463),
            .I(N__19460));
    LocalMux I__1924 (
            .O(N__19460),
            .I(N__19457));
    Span4Mux_h I__1923 (
            .O(N__19457),
            .I(N__19454));
    Span4Mux_v I__1922 (
            .O(N__19454),
            .I(N__19451));
    Odrv4 I__1921 (
            .O(N__19451),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__1920 (
            .O(N__19448),
            .I(N__19445));
    InMux I__1919 (
            .O(N__19445),
            .I(N__19442));
    LocalMux I__1918 (
            .O(N__19442),
            .I(N__19439));
    Span4Mux_h I__1917 (
            .O(N__19439),
            .I(N__19436));
    Odrv4 I__1916 (
            .O(N__19436),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    InMux I__1915 (
            .O(N__19433),
            .I(N__19430));
    LocalMux I__1914 (
            .O(N__19430),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1913 (
            .O(N__19427),
            .I(bfn_2_12_0_));
    InMux I__1912 (
            .O(N__19424),
            .I(N__19421));
    LocalMux I__1911 (
            .O(N__19421),
            .I(N__19418));
    Span4Mux_v I__1910 (
            .O(N__19418),
            .I(N__19415));
    Odrv4 I__1909 (
            .O(N__19415),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__1908 (
            .O(N__19412),
            .I(N__19409));
    InMux I__1907 (
            .O(N__19409),
            .I(N__19406));
    LocalMux I__1906 (
            .O(N__19406),
            .I(N__19403));
    Span4Mux_h I__1905 (
            .O(N__19403),
            .I(N__19400));
    Odrv4 I__1904 (
            .O(N__19400),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1903 (
            .O(N__19397),
            .I(N__19394));
    LocalMux I__1902 (
            .O(N__19394),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1901 (
            .O(N__19391),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    CascadeMux I__1900 (
            .O(N__19388),
            .I(N__19385));
    InMux I__1899 (
            .O(N__19385),
            .I(N__19382));
    LocalMux I__1898 (
            .O(N__19382),
            .I(N__19379));
    Span4Mux_h I__1897 (
            .O(N__19379),
            .I(N__19376));
    Odrv4 I__1896 (
            .O(N__19376),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1895 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__1894 (
            .O(N__19370),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1893 (
            .O(N__19367),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1892 (
            .O(N__19364),
            .I(N__19361));
    LocalMux I__1891 (
            .O(N__19361),
            .I(N__19358));
    Span4Mux_h I__1890 (
            .O(N__19358),
            .I(N__19355));
    Odrv4 I__1889 (
            .O(N__19355),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1888 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__1887 (
            .O(N__19349),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1886 (
            .O(N__19346),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1885 (
            .O(N__19343),
            .I(N__19340));
    InMux I__1884 (
            .O(N__19340),
            .I(N__19337));
    LocalMux I__1883 (
            .O(N__19337),
            .I(N__19334));
    Span4Mux_v I__1882 (
            .O(N__19334),
            .I(N__19331));
    Odrv4 I__1881 (
            .O(N__19331),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1880 (
            .O(N__19328),
            .I(N__19325));
    LocalMux I__1879 (
            .O(N__19325),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1878 (
            .O(N__19322),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1877 (
            .O(N__19319),
            .I(N__19316));
    LocalMux I__1876 (
            .O(N__19316),
            .I(N__19313));
    Span4Mux_v I__1875 (
            .O(N__19313),
            .I(N__19310));
    Odrv4 I__1874 (
            .O(N__19310),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1873 (
            .O(N__19307),
            .I(N__19304));
    LocalMux I__1872 (
            .O(N__19304),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1871 (
            .O(N__19301),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1870 (
            .O(N__19298),
            .I(N__19295));
    InMux I__1869 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__1868 (
            .O(N__19292),
            .I(N__19289));
    Span4Mux_h I__1867 (
            .O(N__19289),
            .I(N__19286));
    Odrv4 I__1866 (
            .O(N__19286),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1865 (
            .O(N__19283),
            .I(N__19280));
    LocalMux I__1864 (
            .O(N__19280),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1863 (
            .O(N__19277),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1862 (
            .O(N__19274),
            .I(N__19271));
    LocalMux I__1861 (
            .O(N__19271),
            .I(N__19268));
    Span4Mux_h I__1860 (
            .O(N__19268),
            .I(N__19265));
    Odrv4 I__1859 (
            .O(N__19265),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1858 (
            .O(N__19262),
            .I(N__19259));
    InMux I__1857 (
            .O(N__19259),
            .I(N__19256));
    LocalMux I__1856 (
            .O(N__19256),
            .I(N__19253));
    Span4Mux_h I__1855 (
            .O(N__19253),
            .I(N__19250));
    Span4Mux_v I__1854 (
            .O(N__19250),
            .I(N__19247));
    Odrv4 I__1853 (
            .O(N__19247),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1852 (
            .O(N__19244),
            .I(N__19241));
    LocalMux I__1851 (
            .O(N__19241),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1850 (
            .O(N__19238),
            .I(N__19235));
    LocalMux I__1849 (
            .O(N__19235),
            .I(N__19232));
    Span4Mux_v I__1848 (
            .O(N__19232),
            .I(N__19229));
    Odrv4 I__1847 (
            .O(N__19229),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1846 (
            .O(N__19226),
            .I(N__19223));
    InMux I__1845 (
            .O(N__19223),
            .I(N__19220));
    LocalMux I__1844 (
            .O(N__19220),
            .I(N__19217));
    Span4Mux_h I__1843 (
            .O(N__19217),
            .I(N__19214));
    Odrv4 I__1842 (
            .O(N__19214),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1841 (
            .O(N__19211),
            .I(N__19208));
    InMux I__1840 (
            .O(N__19208),
            .I(N__19205));
    LocalMux I__1839 (
            .O(N__19205),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1838 (
            .O(N__19202),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1837 (
            .O(N__19199),
            .I(N__19196));
    LocalMux I__1836 (
            .O(N__19196),
            .I(N__19193));
    Span4Mux_v I__1835 (
            .O(N__19193),
            .I(N__19190));
    Odrv4 I__1834 (
            .O(N__19190),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    CascadeMux I__1833 (
            .O(N__19187),
            .I(N__19184));
    InMux I__1832 (
            .O(N__19184),
            .I(N__19181));
    LocalMux I__1831 (
            .O(N__19181),
            .I(N__19178));
    Span4Mux_h I__1830 (
            .O(N__19178),
            .I(N__19175));
    Odrv4 I__1829 (
            .O(N__19175),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    InMux I__1828 (
            .O(N__19172),
            .I(N__19169));
    LocalMux I__1827 (
            .O(N__19169),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1826 (
            .O(N__19166),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1825 (
            .O(N__19163),
            .I(N__19160));
    LocalMux I__1824 (
            .O(N__19160),
            .I(N__19157));
    Span4Mux_s3_h I__1823 (
            .O(N__19157),
            .I(N__19154));
    Span4Mux_v I__1822 (
            .O(N__19154),
            .I(N__19151));
    Odrv4 I__1821 (
            .O(N__19151),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1820 (
            .O(N__19148),
            .I(N__19145));
    InMux I__1819 (
            .O(N__19145),
            .I(N__19142));
    LocalMux I__1818 (
            .O(N__19142),
            .I(N__19139));
    Span4Mux_h I__1817 (
            .O(N__19139),
            .I(N__19136));
    Odrv4 I__1816 (
            .O(N__19136),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    InMux I__1815 (
            .O(N__19133),
            .I(N__19130));
    LocalMux I__1814 (
            .O(N__19130),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1813 (
            .O(N__19127),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1812 (
            .O(N__19124),
            .I(N__19121));
    LocalMux I__1811 (
            .O(N__19121),
            .I(N__19118));
    Span4Mux_v I__1810 (
            .O(N__19118),
            .I(N__19115));
    Odrv4 I__1809 (
            .O(N__19115),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1808 (
            .O(N__19112),
            .I(N__19109));
    InMux I__1807 (
            .O(N__19109),
            .I(N__19106));
    LocalMux I__1806 (
            .O(N__19106),
            .I(N__19103));
    Span4Mux_v I__1805 (
            .O(N__19103),
            .I(N__19100));
    Odrv4 I__1804 (
            .O(N__19100),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1803 (
            .O(N__19097),
            .I(N__19094));
    LocalMux I__1802 (
            .O(N__19094),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1801 (
            .O(N__19091),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1800 (
            .O(N__19088),
            .I(N__19085));
    LocalMux I__1799 (
            .O(N__19085),
            .I(N__19082));
    Span4Mux_v I__1798 (
            .O(N__19082),
            .I(N__19079));
    Odrv4 I__1797 (
            .O(N__19079),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__1796 (
            .O(N__19076),
            .I(N__19073));
    InMux I__1795 (
            .O(N__19073),
            .I(N__19070));
    LocalMux I__1794 (
            .O(N__19070),
            .I(N__19067));
    Span4Mux_v I__1793 (
            .O(N__19067),
            .I(N__19064));
    Odrv4 I__1792 (
            .O(N__19064),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    InMux I__1791 (
            .O(N__19061),
            .I(N__19058));
    LocalMux I__1790 (
            .O(N__19058),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1789 (
            .O(N__19055),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1788 (
            .O(N__19052),
            .I(N__19049));
    LocalMux I__1787 (
            .O(N__19049),
            .I(N__19046));
    Span4Mux_v I__1786 (
            .O(N__19046),
            .I(N__19043));
    Odrv4 I__1785 (
            .O(N__19043),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__1784 (
            .O(N__19040),
            .I(N__19037));
    InMux I__1783 (
            .O(N__19037),
            .I(N__19034));
    LocalMux I__1782 (
            .O(N__19034),
            .I(N__19031));
    Span4Mux_h I__1781 (
            .O(N__19031),
            .I(N__19028));
    Odrv4 I__1780 (
            .O(N__19028),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__1779 (
            .O(N__19025),
            .I(N__19022));
    LocalMux I__1778 (
            .O(N__19022),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1777 (
            .O(N__19019),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1776 (
            .O(N__19016),
            .I(N__19010));
    InMux I__1775 (
            .O(N__19015),
            .I(N__19010));
    LocalMux I__1774 (
            .O(N__19010),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    InMux I__1773 (
            .O(N__19007),
            .I(N__19004));
    LocalMux I__1772 (
            .O(N__19004),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    CascadeMux I__1771 (
            .O(N__19001),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ));
    InMux I__1770 (
            .O(N__18998),
            .I(N__18994));
    InMux I__1769 (
            .O(N__18997),
            .I(N__18991));
    LocalMux I__1768 (
            .O(N__18994),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__1767 (
            .O(N__18991),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__1766 (
            .O(N__18986),
            .I(N__18980));
    InMux I__1765 (
            .O(N__18985),
            .I(N__18980));
    LocalMux I__1764 (
            .O(N__18980),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    InMux I__1763 (
            .O(N__18977),
            .I(N__18974));
    LocalMux I__1762 (
            .O(N__18974),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    CascadeMux I__1761 (
            .O(N__18971),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ));
    CascadeMux I__1760 (
            .O(N__18968),
            .I(N__18964));
    InMux I__1759 (
            .O(N__18967),
            .I(N__18961));
    InMux I__1758 (
            .O(N__18964),
            .I(N__18958));
    LocalMux I__1757 (
            .O(N__18961),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__1756 (
            .O(N__18958),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__1755 (
            .O(N__18953),
            .I(N__18947));
    InMux I__1754 (
            .O(N__18952),
            .I(N__18947));
    LocalMux I__1753 (
            .O(N__18947),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__1752 (
            .O(N__18944),
            .I(N__18941));
    LocalMux I__1751 (
            .O(N__18941),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    CascadeMux I__1750 (
            .O(N__18938),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    InMux I__1749 (
            .O(N__18935),
            .I(N__18932));
    LocalMux I__1748 (
            .O(N__18932),
            .I(N__18928));
    InMux I__1747 (
            .O(N__18931),
            .I(N__18925));
    Odrv4 I__1746 (
            .O(N__18928),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__1745 (
            .O(N__18925),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    CascadeMux I__1744 (
            .O(N__18920),
            .I(N__18917));
    InMux I__1743 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__1742 (
            .O(N__18914),
            .I(N__18911));
    Span4Mux_h I__1741 (
            .O(N__18911),
            .I(N__18906));
    InMux I__1740 (
            .O(N__18910),
            .I(N__18901));
    InMux I__1739 (
            .O(N__18909),
            .I(N__18901));
    Odrv4 I__1738 (
            .O(N__18906),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__1737 (
            .O(N__18901),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__1736 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__1735 (
            .O(N__18893),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    CascadeMux I__1734 (
            .O(N__18890),
            .I(N__18886));
    InMux I__1733 (
            .O(N__18889),
            .I(N__18883));
    InMux I__1732 (
            .O(N__18886),
            .I(N__18880));
    LocalMux I__1731 (
            .O(N__18883),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__1730 (
            .O(N__18880),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    InMux I__1729 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__1728 (
            .O(N__18872),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__1727 (
            .O(N__18869),
            .I(N__18863));
    InMux I__1726 (
            .O(N__18868),
            .I(N__18863));
    LocalMux I__1725 (
            .O(N__18863),
            .I(N__18860));
    Span4Mux_v I__1724 (
            .O(N__18860),
            .I(N__18857));
    Odrv4 I__1723 (
            .O(N__18857),
            .I(\pwm_generator_inst.O_10 ));
    CascadeMux I__1722 (
            .O(N__18854),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ));
    InMux I__1721 (
            .O(N__18851),
            .I(N__18847));
    InMux I__1720 (
            .O(N__18850),
            .I(N__18844));
    LocalMux I__1719 (
            .O(N__18847),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    LocalMux I__1718 (
            .O(N__18844),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__1717 (
            .O(N__18839),
            .I(N__18834));
    InMux I__1716 (
            .O(N__18838),
            .I(N__18831));
    InMux I__1715 (
            .O(N__18837),
            .I(N__18828));
    LocalMux I__1714 (
            .O(N__18834),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__1713 (
            .O(N__18831),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__1712 (
            .O(N__18828),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    CascadeMux I__1711 (
            .O(N__18821),
            .I(N__18818));
    InMux I__1710 (
            .O(N__18818),
            .I(N__18815));
    LocalMux I__1709 (
            .O(N__18815),
            .I(N__18812));
    Odrv4 I__1708 (
            .O(N__18812),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    CascadeMux I__1707 (
            .O(N__18809),
            .I(N__18805));
    InMux I__1706 (
            .O(N__18808),
            .I(N__18802));
    InMux I__1705 (
            .O(N__18805),
            .I(N__18799));
    LocalMux I__1704 (
            .O(N__18802),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1703 (
            .O(N__18799),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    CascadeMux I__1702 (
            .O(N__18794),
            .I(N__18791));
    InMux I__1701 (
            .O(N__18791),
            .I(N__18785));
    InMux I__1700 (
            .O(N__18790),
            .I(N__18785));
    LocalMux I__1699 (
            .O(N__18785),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1698 (
            .O(N__18782),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__1697 (
            .O(N__18779),
            .I(N__18776));
    LocalMux I__1696 (
            .O(N__18776),
            .I(N__18771));
    InMux I__1695 (
            .O(N__18775),
            .I(N__18766));
    InMux I__1694 (
            .O(N__18774),
            .I(N__18766));
    Span4Mux_s1_h I__1693 (
            .O(N__18771),
            .I(N__18763));
    LocalMux I__1692 (
            .O(N__18766),
            .I(pwm_duty_input_7));
    Odrv4 I__1691 (
            .O(N__18763),
            .I(pwm_duty_input_7));
    InMux I__1690 (
            .O(N__18758),
            .I(N__18753));
    InMux I__1689 (
            .O(N__18757),
            .I(N__18748));
    InMux I__1688 (
            .O(N__18756),
            .I(N__18748));
    LocalMux I__1687 (
            .O(N__18753),
            .I(N__18745));
    LocalMux I__1686 (
            .O(N__18748),
            .I(pwm_duty_input_5));
    Odrv4 I__1685 (
            .O(N__18745),
            .I(pwm_duty_input_5));
    InMux I__1684 (
            .O(N__18740),
            .I(N__18736));
    CascadeMux I__1683 (
            .O(N__18739),
            .I(N__18733));
    LocalMux I__1682 (
            .O(N__18736),
            .I(N__18729));
    InMux I__1681 (
            .O(N__18733),
            .I(N__18724));
    InMux I__1680 (
            .O(N__18732),
            .I(N__18724));
    Span4Mux_s2_h I__1679 (
            .O(N__18729),
            .I(N__18721));
    LocalMux I__1678 (
            .O(N__18724),
            .I(pwm_duty_input_8));
    Odrv4 I__1677 (
            .O(N__18721),
            .I(pwm_duty_input_8));
    InMux I__1676 (
            .O(N__18716),
            .I(N__18713));
    LocalMux I__1675 (
            .O(N__18713),
            .I(N__18708));
    InMux I__1674 (
            .O(N__18712),
            .I(N__18703));
    InMux I__1673 (
            .O(N__18711),
            .I(N__18703));
    Span4Mux_s2_h I__1672 (
            .O(N__18708),
            .I(N__18700));
    LocalMux I__1671 (
            .O(N__18703),
            .I(pwm_duty_input_9));
    Odrv4 I__1670 (
            .O(N__18700),
            .I(pwm_duty_input_9));
    CascadeMux I__1669 (
            .O(N__18695),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__1668 (
            .O(N__18692),
            .I(N__18687));
    InMux I__1667 (
            .O(N__18691),
            .I(N__18682));
    InMux I__1666 (
            .O(N__18690),
            .I(N__18682));
    LocalMux I__1665 (
            .O(N__18687),
            .I(N__18679));
    LocalMux I__1664 (
            .O(N__18682),
            .I(N__18676));
    Span4Mux_s1_h I__1663 (
            .O(N__18679),
            .I(N__18673));
    Odrv4 I__1662 (
            .O(N__18676),
            .I(pwm_duty_input_6));
    Odrv4 I__1661 (
            .O(N__18673),
            .I(pwm_duty_input_6));
    InMux I__1660 (
            .O(N__18668),
            .I(N__18659));
    InMux I__1659 (
            .O(N__18667),
            .I(N__18659));
    InMux I__1658 (
            .O(N__18666),
            .I(N__18659));
    LocalMux I__1657 (
            .O(N__18659),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1656 (
            .O(N__18656),
            .I(N__18652));
    InMux I__1655 (
            .O(N__18655),
            .I(N__18649));
    LocalMux I__1654 (
            .O(N__18652),
            .I(pwm_duty_input_0));
    LocalMux I__1653 (
            .O(N__18649),
            .I(pwm_duty_input_0));
    InMux I__1652 (
            .O(N__18644),
            .I(N__18640));
    InMux I__1651 (
            .O(N__18643),
            .I(N__18637));
    LocalMux I__1650 (
            .O(N__18640),
            .I(pwm_duty_input_2));
    LocalMux I__1649 (
            .O(N__18637),
            .I(pwm_duty_input_2));
    InMux I__1648 (
            .O(N__18632),
            .I(N__18628));
    InMux I__1647 (
            .O(N__18631),
            .I(N__18625));
    LocalMux I__1646 (
            .O(N__18628),
            .I(pwm_duty_input_1));
    LocalMux I__1645 (
            .O(N__18625),
            .I(pwm_duty_input_1));
    InMux I__1644 (
            .O(N__18620),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1643 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__1642 (
            .O(N__18614),
            .I(N__18610));
    InMux I__1641 (
            .O(N__18613),
            .I(N__18607));
    Odrv4 I__1640 (
            .O(N__18610),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1639 (
            .O(N__18607),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    CascadeMux I__1638 (
            .O(N__18602),
            .I(N__18599));
    InMux I__1637 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__1636 (
            .O(N__18596),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1635 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__1634 (
            .O(N__18590),
            .I(un7_start_stop_0_a3));
    InMux I__1633 (
            .O(N__18587),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__1632 (
            .O(N__18584),
            .I(bfn_1_11_0_));
    InMux I__1631 (
            .O(N__18581),
            .I(N__18577));
    InMux I__1630 (
            .O(N__18580),
            .I(N__18574));
    LocalMux I__1629 (
            .O(N__18577),
            .I(N__18569));
    LocalMux I__1628 (
            .O(N__18574),
            .I(N__18569));
    Span4Mux_v I__1627 (
            .O(N__18569),
            .I(N__18566));
    Odrv4 I__1626 (
            .O(N__18566),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1625 (
            .O(N__18563),
            .I(N__18560));
    LocalMux I__1624 (
            .O(N__18560),
            .I(N__18557));
    Span4Mux_v I__1623 (
            .O(N__18557),
            .I(N__18554));
    Odrv4 I__1622 (
            .O(N__18554),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1621 (
            .O(N__18551),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1620 (
            .O(N__18548),
            .I(N__18545));
    LocalMux I__1619 (
            .O(N__18545),
            .I(N__18542));
    Span4Mux_v I__1618 (
            .O(N__18542),
            .I(N__18539));
    Odrv4 I__1617 (
            .O(N__18539),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1616 (
            .O(N__18536),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1615 (
            .O(N__18533),
            .I(N__18530));
    LocalMux I__1614 (
            .O(N__18530),
            .I(N__18527));
    Span4Mux_v I__1613 (
            .O(N__18527),
            .I(N__18524));
    Odrv4 I__1612 (
            .O(N__18524),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1611 (
            .O(N__18521),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1610 (
            .O(N__18518),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    InMux I__1609 (
            .O(N__18515),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1608 (
            .O(N__18512),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1607 (
            .O(N__18509),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1606 (
            .O(N__18506),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1605 (
            .O(N__18503),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1604 (
            .O(N__18500),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__1603 (
            .O(N__18497),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__1602 (
            .O(N__18494),
            .I(bfn_1_9_0_));
    InMux I__1601 (
            .O(N__18491),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__1600 (
            .O(N__18488),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__1599 (
            .O(N__18485),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__1598 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__1597 (
            .O(N__18479),
            .I(N__18476));
    Odrv4 I__1596 (
            .O(N__18476),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1595 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__1594 (
            .O(N__18470),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1593 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__1592 (
            .O(N__18464),
            .I(N__18461));
    Span4Mux_h I__1591 (
            .O(N__18461),
            .I(N__18458));
    Odrv4 I__1590 (
            .O(N__18458),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1589 (
            .O(N__18455),
            .I(N__18452));
    LocalMux I__1588 (
            .O(N__18452),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1587 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__1586 (
            .O(N__18446),
            .I(N__18443));
    Odrv4 I__1585 (
            .O(N__18443),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1584 (
            .O(N__18440),
            .I(N__18437));
    LocalMux I__1583 (
            .O(N__18437),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1582 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__1581 (
            .O(N__18431),
            .I(N__18428));
    Span4Mux_h I__1580 (
            .O(N__18428),
            .I(N__18425));
    Odrv4 I__1579 (
            .O(N__18425),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1578 (
            .O(N__18422),
            .I(N__18419));
    LocalMux I__1577 (
            .O(N__18419),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__1576 (
            .O(N__18416),
            .I(N__18413));
    LocalMux I__1575 (
            .O(N__18413),
            .I(N__18410));
    Span4Mux_v I__1574 (
            .O(N__18410),
            .I(N__18407));
    Odrv4 I__1573 (
            .O(N__18407),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1572 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__1571 (
            .O(N__18401),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__1570 (
            .O(N__18398),
            .I(N__18395));
    LocalMux I__1569 (
            .O(N__18395),
            .I(N__18392));
    Odrv4 I__1568 (
            .O(N__18392),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1567 (
            .O(N__18389),
            .I(N__18386));
    LocalMux I__1566 (
            .O(N__18386),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__1565 (
            .O(N__18383),
            .I(N__18380));
    LocalMux I__1564 (
            .O(N__18380),
            .I(N__18377));
    Odrv4 I__1563 (
            .O(N__18377),
            .I(\pwm_generator_inst.O_9 ));
    CascadeMux I__1562 (
            .O(N__18374),
            .I(N__18371));
    InMux I__1561 (
            .O(N__18371),
            .I(N__18368));
    LocalMux I__1560 (
            .O(N__18368),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1559 (
            .O(N__18365),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1558 (
            .O(N__18362),
            .I(N__18359));
    LocalMux I__1557 (
            .O(N__18359),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__1556 (
            .O(N__18356),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    CascadeMux I__1555 (
            .O(N__18353),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_ ));
    InMux I__1554 (
            .O(N__18350),
            .I(N__18344));
    InMux I__1553 (
            .O(N__18349),
            .I(N__18344));
    LocalMux I__1552 (
            .O(N__18344),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1551 (
            .O(N__18341),
            .I(N__18329));
    InMux I__1550 (
            .O(N__18340),
            .I(N__18329));
    InMux I__1549 (
            .O(N__18339),
            .I(N__18329));
    InMux I__1548 (
            .O(N__18338),
            .I(N__18329));
    LocalMux I__1547 (
            .O(N__18329),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__1546 (
            .O(N__18326),
            .I(N__18323));
    LocalMux I__1545 (
            .O(N__18323),
            .I(N__18320));
    Odrv4 I__1544 (
            .O(N__18320),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1543 (
            .O(N__18317),
            .I(N__18314));
    LocalMux I__1542 (
            .O(N__18314),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1541 (
            .O(N__18311),
            .I(N__18308));
    LocalMux I__1540 (
            .O(N__18308),
            .I(N__18305));
    Span4Mux_v I__1539 (
            .O(N__18305),
            .I(N__18302));
    Odrv4 I__1538 (
            .O(N__18302),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1537 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__1536 (
            .O(N__18296),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1535 (
            .O(N__18293),
            .I(N__18290));
    LocalMux I__1534 (
            .O(N__18290),
            .I(N__18287));
    Odrv4 I__1533 (
            .O(N__18287),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1532 (
            .O(N__18284),
            .I(N__18281));
    LocalMux I__1531 (
            .O(N__18281),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    CascadeMux I__1530 (
            .O(N__18278),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    CascadeMux I__1529 (
            .O(N__18275),
            .I(\current_shift_inst.PI_CTRL.N_27_cascade_ ));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_6 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_14 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_22 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_30 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(un5_counter_cry_8),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_8 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_16 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_24 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.z_cry_7 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.z_cry_15 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.z_cry_23 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_8 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_16 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_24 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_7 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_8_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_23_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_15 ),
            .carryinitout(bfn_8_23_0_));
    defparam IN_MUX_bfv_8_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_24_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_23 ),
            .carryinitout(bfn_8_24_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_15 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_23 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryinitout(bfn_11_13_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__34067),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_335_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__24020),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_187_i_g ));
    ICE_GB \current_shift_inst.timer_phase.running_RNIC90O_0  (
            .USERSIGNALTOGLOBALBUFFER(N__27425),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_phase.N_188_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__22857),
            .CLKHFEN(N__22859),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__22858),
            .RGB2PWM(N__19601),
            .RGB1(rgb_g),
            .CURREN(N__22993),
            .RGB2(rgb_b),
            .RGB1PWM(N__18593),
            .RGB0PWM(N__47463),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_4_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_4_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_4_4 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_4_4  (
            .in0(N__21323),
            .in1(N__19892),
            .in2(N__21896),
            .in3(N__19829),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48008),
            .ce(N__32559),
            .sr(N__47350));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_1_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_1_5_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__21208),
            .in2(_gnd_net_),
            .in3(N__21349),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_5_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_5_1  (
            .in0(N__21247),
            .in1(N__21286),
            .in2(N__18278),
            .in3(N__21322),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(\current_shift_inst.PI_CTRL.N_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_2 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_2  (
            .in0(N__19828),
            .in1(N__20870),
            .in2(N__18275),
            .in3(N__19589),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48007),
            .ce(N__32560),
            .sr(N__47357));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_3 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_3  (
            .in0(N__21350),
            .in1(N__19890),
            .in2(N__21893),
            .in3(N__19826),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48007),
            .ce(N__32560),
            .sr(N__47357));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_5 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_5  (
            .in0(N__21287),
            .in1(N__19891),
            .in2(N__21894),
            .in3(N__19827),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48007),
            .ce(N__32560),
            .sr(N__47357));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_0  (
            .in0(N__18668),
            .in1(N__18340),
            .in2(N__20930),
            .in3(N__18350),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48005),
            .ce(N__32540),
            .sr(N__47367));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_6_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_6_1  (
            .in0(N__20990),
            .in1(N__18362),
            .in2(N__21895),
            .in3(N__19813),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_6_2 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_6_2  (
            .in0(N__19886),
            .in1(N__20896),
            .in2(N__18356),
            .in3(N__18790),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3  (
            .in0(N__18339),
            .in1(N__20945),
            .in2(N__18353),
            .in3(N__18667),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48005),
            .ce(N__32540),
            .sr(N__47367));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_4  (
            .in0(N__18666),
            .in1(N__18338),
            .in2(N__20963),
            .in3(N__18349),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48005),
            .ce(N__32540),
            .sr(N__47367));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_5 .LUT_INIT=16'b1101110111001101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_5  (
            .in0(N__18341),
            .in1(N__20897),
            .in2(N__18794),
            .in3(N__19887),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48005),
            .ce(N__32540),
            .sr(N__47367));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0  (
            .in0(N__18326),
            .in1(N__18317),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__18299),
            .in2(_gnd_net_),
            .in3(N__18311),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__18284),
            .in2(_gnd_net_),
            .in3(N__18293),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__18473),
            .in2(_gnd_net_),
            .in3(N__18482),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__18455),
            .in2(_gnd_net_),
            .in3(N__18467),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__18440),
            .in2(_gnd_net_),
            .in3(N__18449),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__18422),
            .in2(_gnd_net_),
            .in3(N__18434),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(N__18404),
            .in2(_gnd_net_),
            .in3(N__18416),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0  (
            .in0(N__18398),
            .in1(N__18389),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18374),
            .in3(N__18383),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18890),
            .in3(N__18365),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3  (
            .in0(N__20030),
            .in1(N__18581),
            .in2(_gnd_net_),
            .in3(N__18509),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__20098),
            .in2(_gnd_net_),
            .in3(N__18506),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__20163),
            .in2(_gnd_net_),
            .in3(N__18503),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__18837),
            .in2(_gnd_net_),
            .in3(N__18500),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18809),
            .in3(N__18497),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__18997),
            .in2(_gnd_net_),
            .in3(N__18494),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18968),
            .in3(N__18491),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__18909),
            .in2(_gnd_net_),
            .in3(N__18488),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18485),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__18839),
            .in2(_gnd_net_),
            .in3(N__18850),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_7  (
            .in0(N__18910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18931),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__18580),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__18563),
            .in2(_gnd_net_),
            .in3(N__18551),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__18548),
            .in2(_gnd_net_),
            .in3(N__18536),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18533),
            .in2(_gnd_net_),
            .in3(N__18521),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__19244),
            .in2(_gnd_net_),
            .in3(N__18518),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__22994),
            .in2(N__19211),
            .in3(N__18515),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__19172),
            .in2(N__23055),
            .in3(N__18512),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__19133),
            .in2(N__23056),
            .in3(N__18587),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__19097),
            .in2(_gnd_net_),
            .in3(N__18584),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__19061),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__19025),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__19472),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__19433),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__19397),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__19373),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__19352),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__19328),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__19307),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__19283),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__19625),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18620),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5  (
            .in0(N__18613),
            .in1(N__19672),
            .in2(_gnd_net_),
            .in3(N__20615),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_0 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_0  (
            .in0(N__19676),
            .in1(N__18617),
            .in2(N__18602),
            .in3(N__20614),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_1_29_0 .C_ON=1'b0;
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_1_29_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \current_shift_inst.un7_start_stop_0_a3_LC_1_29_0  (
            .in0(N__47462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33731),
            .lcout(un7_start_stop_0_a3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_2_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_2_5_0 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_2_5_0  (
            .in0(N__21248),
            .in1(N__19888),
            .in2(N__21891),
            .in3(N__19814),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48006),
            .ce(N__32548),
            .sr(N__47351));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_2_5_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_2_5_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_2_5_6 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_2_5_6  (
            .in0(N__21209),
            .in1(N__19889),
            .in2(N__21892),
            .in3(N__19815),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48006),
            .ce(N__32548),
            .sr(N__47351));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_0 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_0  (
            .in0(N__19575),
            .in1(N__21861),
            .in2(_gnd_net_),
            .in3(N__20859),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_1  (
            .in0(N__18775),
            .in1(N__18712),
            .in2(N__18739),
            .in3(N__18691),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_2  (
            .in0(N__19555),
            .in1(N__19518),
            .in2(N__18782),
            .in3(N__18757),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__18774),
            .in2(_gnd_net_),
            .in3(N__18756),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_5  (
            .in0(N__18732),
            .in1(N__18711),
            .in2(N__18695),
            .in3(N__18690),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_6_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_6_6  (
            .in0(N__19576),
            .in1(N__21862),
            .in2(_gnd_net_),
            .in3(N__19885),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_6_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_6_7  (
            .in0(N__18656),
            .in1(N__18644),
            .in2(_gnd_net_),
            .in3(N__18632),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_7_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_7_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_7_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_2_7_5  (
            .in0(N__20420),
            .in1(N__20360),
            .in2(N__20553),
            .in3(N__19730),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48003),
            .ce(),
            .sr(N__47368));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_2_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_2_7_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_2_7_7  (
            .in0(N__20421),
            .in1(N__20361),
            .in2(N__20554),
            .in3(N__19721),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48003),
            .ce(),
            .sr(N__47368));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_0 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_0  (
            .in0(N__18935),
            .in1(N__20032),
            .in2(N__18920),
            .in3(N__18896),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_1  (
            .in0(N__18868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18889),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_2 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_2  (
            .in0(N__18875),
            .in1(N__18869),
            .in2(N__18854),
            .in3(N__20031),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_2_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_2_8_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_2_8_4  (
            .in0(N__34990),
            .in1(N__35617),
            .in2(N__40553),
            .in3(N__39596),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48000),
            .ce(N__33569),
            .sr(N__47375));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_2_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_2_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_2_8_5 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_2_8_5  (
            .in0(N__35616),
            .in1(N__36418),
            .in2(N__40559),
            .in3(N__34989),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48000),
            .ce(N__33569),
            .sr(N__47375));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_2_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_2_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_2_8_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_2_8_6  (
            .in0(N__34991),
            .in1(_gnd_net_),
            .in2(N__34691),
            .in3(N__40554),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48000),
            .ce(N__33569),
            .sr(N__47375));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0  (
            .in0(N__18851),
            .in1(N__18838),
            .in2(N__18821),
            .in3(N__20034),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1  (
            .in0(N__18808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19015),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2  (
            .in0(N__19016),
            .in1(N__19007),
            .in2(N__19001),
            .in3(N__20035),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__18985),
            .in2(_gnd_net_),
            .in3(N__18998),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_4  (
            .in0(N__18986),
            .in1(N__18977),
            .in2(N__18971),
            .in3(N__20033),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__18952),
            .in2(_gnd_net_),
            .in3(N__18967),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_6  (
            .in0(N__18953),
            .in1(N__18944),
            .in2(N__18938),
            .in3(N__20036),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__20167),
            .in2(_gnd_net_),
            .in3(N__20140),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_2_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_2_10_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_2_10_0 .LUT_INIT=16'b1111010111110011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_2_10_0  (
            .in0(N__20430),
            .in1(N__20401),
            .in2(N__19940),
            .in3(N__20597),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47996),
            .ce(),
            .sr(N__47388));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_10_2 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_2_10_2  (
            .in0(N__20431),
            .in1(N__20402),
            .in2(N__19901),
            .in3(N__20598),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47996),
            .ce(),
            .sr(N__47388));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_10_3  (
            .in0(N__20068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20097),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__19274),
            .in2(N__19262),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__19238),
            .in2(N__19226),
            .in3(N__19202),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__19199),
            .in2(N__19187),
            .in3(N__19166),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__19163),
            .in2(N__19148),
            .in3(N__19127),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__19124),
            .in2(N__19112),
            .in3(N__19091),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__19088),
            .in2(N__19076),
            .in3(N__19055),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__19052),
            .in2(N__19040),
            .in3(N__19019),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__19499),
            .in2(N__19487),
            .in3(N__19466),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__19463),
            .in2(N__19448),
            .in3(N__19427),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__19424),
            .in2(N__19412),
            .in3(N__19391),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__19657),
            .in2(N__19388),
            .in3(N__19367),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__19364),
            .in2(N__19673),
            .in3(N__19346),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__19661),
            .in2(N__19343),
            .in3(N__19322),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__19319),
            .in2(N__19674),
            .in3(N__19301),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__19665),
            .in2(N__19298),
            .in3(N__19277),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__19682),
            .in2(N__19675),
            .in3(N__19619),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0  (
            .in0(N__19616),
            .in1(N__19610),
            .in2(_gnd_net_),
            .in3(N__19604),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.N_32_i_i_LC_2_29_5 .C_ON=1'b0;
    defparam \current_shift_inst.N_32_i_i_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.N_32_i_i_LC_2_29_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.N_32_i_i_LC_2_29_5  (
            .in0(_gnd_net_),
            .in1(N__33730),
            .in2(_gnd_net_),
            .in3(N__47461),
            .lcout(N_32_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_1 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_1  (
            .in0(N__20866),
            .in1(N__19577),
            .in2(N__21890),
            .in3(N__19863),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_0_5_LC_3_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_0_5_LC_3_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_0_5_LC_3_6_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_0_5_LC_3_6_1  (
            .in0(_gnd_net_),
            .in1(N__21201),
            .in2(_gnd_net_),
            .in3(N__21343),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_3_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_3_6_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_3_6_2  (
            .in0(N__21240),
            .in1(N__21279),
            .in2(N__19580),
            .in3(N__21315),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_6 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_6  (
            .in0(N__19562),
            .in1(N__19556),
            .in2(N__19535),
            .in3(N__19526),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_3_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_3_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_3_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_3_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21860),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48001),
            .ce(N__32547),
            .sr(N__47358));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_3_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27836),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48001),
            .ce(N__32547),
            .sr(N__47358));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_3_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_3_7_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_3_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_3_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27965),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48001),
            .ce(N__32547),
            .sr(N__47358));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0  (
            .in0(_gnd_net_),
            .in1(N__19751),
            .in2(N__20042),
            .in3(N__20041),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19745),
            .in3(N__19733),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(N__19967),
            .in2(_gnd_net_),
            .in3(N__19724),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(N__20111),
            .in2(_gnd_net_),
            .in3(N__19715),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(N__19712),
            .in2(_gnd_net_),
            .in3(N__19706),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(N__19703),
            .in2(_gnd_net_),
            .in3(N__19697),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6  (
            .in0(_gnd_net_),
            .in1(N__19694),
            .in2(_gnd_net_),
            .in3(N__19685),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7  (
            .in0(_gnd_net_),
            .in1(N__19958),
            .in2(_gnd_net_),
            .in3(N__19952),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19949),
            .in3(N__19931),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1  (
            .in0(N__19928),
            .in1(N__20040),
            .in2(N__19919),
            .in3(N__19904),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_3_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_3_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_3_9_6  (
            .in0(N__19775),
            .in1(N__20189),
            .in2(N__19760),
            .in3(N__20333),
            .lcout(\current_shift_inst.PI_CTRL.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_9_7  (
            .in0(N__20651),
            .in1(N__20204),
            .in2(N__20180),
            .in3(N__19766),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINKF4_12_LC_3_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINKF4_12_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINKF4_12_LC_3_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINKF4_12_LC_3_10_0  (
            .in0(N__21557),
            .in1(N__21107),
            .in2(N__21932),
            .in3(N__21575),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRO62_11_LC_3_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRO62_11_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRO62_11_LC_3_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRO62_11_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__21556),
            .in2(_gnd_net_),
            .in3(N__21137),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4TS8_10_LC_3_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4TS8_10_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4TS8_10_LC_3_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4TS8_10_LC_3_10_2  (
            .in0(N__21160),
            .in1(N__20198),
            .in2(N__19769),
            .in3(N__21574),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID6B4_10_LC_3_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID6B4_10_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID6B4_10_LC_3_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNID6B4_10_LC_3_10_3  (
            .in0(N__21515),
            .in1(N__21473),
            .in2(N__21539),
            .in3(N__21161),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_20_LC_3_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_20_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_20_LC_3_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_20_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(N__21664),
            .in2(_gnd_net_),
            .in3(N__21383),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIR5H5_12_LC_3_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIR5H5_12_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIR5H5_12_LC_3_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIR5H5_12_LC_3_10_6  (
            .in0(N__21625),
            .in1(N__21514),
            .in2(N__20207),
            .in3(N__21106),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_19_LC_3_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_19_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_19_LC_3_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_19_LC_3_11_1  (
            .in0(N__21701),
            .in1(N__21719),
            .in2(N__21931),
            .in3(N__21406),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1U52_18_LC_3_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1U52_18_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1U52_18_LC_3_11_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1U52_18_LC_3_11_4  (
            .in0(N__21407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21425),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_20_LC_3_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_20_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_20_LC_3_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_20_LC_3_11_5  (
            .in0(N__21644),
            .in1(N__21382),
            .in2(N__20192),
            .in3(N__21595),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINID4_13_LC_3_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINID4_13_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINID4_13_LC_3_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINID4_13_LC_3_11_6  (
            .in0(N__21469),
            .in1(N__21643),
            .in2(N__21596),
            .in3(N__21538),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_3_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_3_12_1 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_3_12_1  (
            .in0(N__20168),
            .in1(N__20147),
            .in2(N__20129),
            .in3(N__19996),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_12_5 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_12_5  (
            .in0(N__20099),
            .in1(N__20075),
            .in2(N__20057),
            .in3(N__19995),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_counter_cry_1_c_LC_4_5_0.C_ON=1'b1;
    defparam un5_counter_cry_1_c_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam un5_counter_cry_1_c_LC_4_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_counter_cry_1_c_LC_4_5_0 (
            .in0(_gnd_net_),
            .in1(N__20704),
            .in2(N__20686),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(un5_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_4_5_1.C_ON=1'b1;
    defparam counter_2_LC_4_5_1.SEQ_MODE=4'b1010;
    defparam counter_2_LC_4_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_2_LC_4_5_1 (
            .in0(_gnd_net_),
            .in1(N__20269),
            .in2(_gnd_net_),
            .in3(N__20231),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(un5_counter_cry_1),
            .carryout(un5_counter_cry_2),
            .clk(N__48004),
            .ce(),
            .sr(N__47328));
    defparam counter_3_LC_4_5_2.C_ON=1'b1;
    defparam counter_3_LC_4_5_2.SEQ_MODE=4'b1010;
    defparam counter_3_LC_4_5_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_3_LC_4_5_2 (
            .in0(_gnd_net_),
            .in1(N__20792),
            .in2(_gnd_net_),
            .in3(N__20228),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(un5_counter_cry_2),
            .carryout(un5_counter_cry_3),
            .clk(N__48004),
            .ce(),
            .sr(N__47328));
    defparam counter_4_LC_4_5_3.C_ON=1'b1;
    defparam counter_4_LC_4_5_3.SEQ_MODE=4'b1010;
    defparam counter_4_LC_4_5_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_4_LC_4_5_3 (
            .in0(_gnd_net_),
            .in1(N__20804),
            .in2(_gnd_net_),
            .in3(N__20225),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(un5_counter_cry_3),
            .carryout(un5_counter_cry_4),
            .clk(N__48004),
            .ce(),
            .sr(N__47328));
    defparam counter_5_LC_4_5_4.C_ON=1'b1;
    defparam counter_5_LC_4_5_4.SEQ_MODE=4'b1010;
    defparam counter_5_LC_4_5_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_5_LC_4_5_4 (
            .in0(_gnd_net_),
            .in1(N__20780),
            .in2(_gnd_net_),
            .in3(N__20222),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(un5_counter_cry_4),
            .carryout(un5_counter_cry_5),
            .clk(N__48004),
            .ce(),
            .sr(N__47328));
    defparam counter_6_LC_4_5_5.C_ON=1'b1;
    defparam counter_6_LC_4_5_5.SEQ_MODE=4'b1010;
    defparam counter_6_LC_4_5_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_6_LC_4_5_5 (
            .in0(_gnd_net_),
            .in1(N__20768),
            .in2(_gnd_net_),
            .in3(N__20219),
            .lcout(counterZ0Z_6),
            .ltout(),
            .carryin(un5_counter_cry_5),
            .carryout(un5_counter_cry_6),
            .clk(N__48004),
            .ce(),
            .sr(N__47328));
    defparam counter_RNO_0_7_LC_4_5_6.C_ON=1'b1;
    defparam counter_RNO_0_7_LC_4_5_6.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_7_LC_4_5_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_7_LC_4_5_6 (
            .in0(_gnd_net_),
            .in1(N__20630),
            .in2(_gnd_net_),
            .in3(N__20216),
            .lcout(counter_RNO_0Z0Z_7),
            .ltout(),
            .carryin(un5_counter_cry_6),
            .carryout(un5_counter_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_8_LC_4_5_7.C_ON=1'b1;
    defparam counter_8_LC_4_5_7.SEQ_MODE=4'b1010;
    defparam counter_8_LC_4_5_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_8_LC_4_5_7 (
            .in0(_gnd_net_),
            .in1(N__20284),
            .in2(_gnd_net_),
            .in3(N__20213),
            .lcout(counterZ0Z_8),
            .ltout(),
            .carryin(un5_counter_cry_7),
            .carryout(un5_counter_cry_8),
            .clk(N__48004),
            .ce(),
            .sr(N__47328));
    defparam counter_9_LC_4_6_0.C_ON=1'b1;
    defparam counter_9_LC_4_6_0.SEQ_MODE=4'b1010;
    defparam counter_9_LC_4_6_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_9_LC_4_6_0 (
            .in0(_gnd_net_),
            .in1(N__20297),
            .in2(_gnd_net_),
            .in3(N__20210),
            .lcout(counterZ0Z_9),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(un5_counter_cry_9),
            .clk(N__48002),
            .ce(),
            .sr(N__47341));
    defparam counter_RNO_0_10_LC_4_6_1.C_ON=1'b1;
    defparam counter_RNO_0_10_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_10_LC_4_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_10_LC_4_6_1 (
            .in0(_gnd_net_),
            .in1(N__20719),
            .in2(_gnd_net_),
            .in3(N__20321),
            .lcout(counter_RNO_0Z0Z_10),
            .ltout(),
            .carryin(un5_counter_cry_9),
            .carryout(un5_counter_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_11_LC_4_6_2.C_ON=1'b1;
    defparam counter_11_LC_4_6_2.SEQ_MODE=4'b1010;
    defparam counter_11_LC_4_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_11_LC_4_6_2 (
            .in0(_gnd_net_),
            .in1(N__20311),
            .in2(_gnd_net_),
            .in3(N__20318),
            .lcout(counterZ0Z_11),
            .ltout(),
            .carryin(un5_counter_cry_10),
            .carryout(un5_counter_cry_11),
            .clk(N__48002),
            .ce(),
            .sr(N__47341));
    defparam counter_RNO_0_12_LC_4_6_3.C_ON=1'b0;
    defparam counter_RNO_0_12_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_12_LC_4_6_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_RNO_0_12_LC_4_6_3 (
            .in0(_gnd_net_),
            .in1(N__20743),
            .in2(_gnd_net_),
            .in3(N__20315),
            .lcout(counter_RNO_0Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIM6001_12_LC_4_7_0.C_ON=1'b0;
    defparam counter_RNIM6001_12_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam counter_RNIM6001_12_LC_4_7_0.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNIM6001_12_LC_4_7_0 (
            .in0(N__20312),
            .in1(N__20296),
            .in2(N__20744),
            .in3(N__20285),
            .lcout(un2_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIRTIM_1_LC_4_7_3.C_ON=1'b0;
    defparam counter_RNIRTIM_1_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam counter_RNIRTIM_1_LC_4_7_3.LUT_INIT=16'b0000000001000000;
    LogicCell40 counter_RNIRTIM_1_LC_4_7_3 (
            .in0(N__20270),
            .in1(N__20626),
            .in2(N__20720),
            .in3(N__20703),
            .lcout(un2_counter_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_0 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_4_8_0  (
            .in0(N__20513),
            .in1(N__20447),
            .in2(N__20397),
            .in3(N__20255),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_8_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_8_1 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_4_8_1  (
            .in0(N__20446),
            .in1(N__20379),
            .in2(N__20556),
            .in3(N__20249),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_8_2 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_4_8_2  (
            .in0(N__20514),
            .in1(N__20448),
            .in2(N__20398),
            .in3(N__20243),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_8_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_8_3 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_4_8_3  (
            .in0(N__20445),
            .in1(N__20237),
            .in2(N__20555),
            .in3(N__20378),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_8_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_8_4 .LUT_INIT=16'b1111111100100111;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_4_8_4  (
            .in0(N__20515),
            .in1(N__20449),
            .in2(N__20399),
            .in3(N__20645),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam counter_7_LC_4_8_5.C_ON=1'b0;
    defparam counter_7_LC_4_8_5.SEQ_MODE=4'b1010;
    defparam counter_7_LC_4_8_5.LUT_INIT=16'b0100110011001100;
    LogicCell40 counter_7_LC_4_8_5 (
            .in0(N__21056),
            .in1(N__20639),
            .in2(N__21092),
            .in3(N__21026),
            .lcout(counterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_8_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_8_6 .LUT_INIT=16'b1111111100100111;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_4_8_6  (
            .in0(N__20516),
            .in1(N__20450),
            .in2(N__20400),
            .in3(N__20342),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__47359));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28412),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47994),
            .ce(N__32485),
            .sr(N__47369));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27656),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47994),
            .ce(N__32485),
            .sr(N__47369));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28184),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47994),
            .ce(N__32485),
            .sr(N__47369));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_17_LC_4_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_17_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_17_LC_4_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_17_LC_4_10_1  (
            .in0(N__21448),
            .in1(N__21700),
            .in2(N__21626),
            .in3(N__21665),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_11_LC_4_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_11_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_11_LC_4_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_11_LC_4_10_2  (
            .in0(N__21494),
            .in1(N__20327),
            .in2(N__20336),
            .in3(N__21136),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_21_LC_4_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_21_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_21_LC_4_10_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_21_LC_4_10_3  (
            .in0(N__21682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21718),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_4_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_4_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_4_10_5  (
            .in0(N__21683),
            .in1(N__21493),
            .in2(N__21449),
            .in3(N__21424),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28339),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47987),
            .ce(N__32490),
            .sr(N__47381));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_4_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_4_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_4_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28876),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47987),
            .ce(N__32490),
            .sr(N__47381));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_4_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28792),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47987),
            .ce(N__32490),
            .sr(N__47381));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_4_11_6  (
            .in0(N__28108),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47987),
            .ce(N__32490),
            .sr(N__47381));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29447),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47987),
            .ce(N__32490),
            .sr(N__47381));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28030),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__32497),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_4_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_4_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_4_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29335),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__32497),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29146),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__32497),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28633),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__32497),
            .sr(N__47389));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_6 (
            .in0(N__20831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIN1J6_3_LC_5_5_2.C_ON=1'b0;
    defparam counter_RNIN1J6_3_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam counter_RNIN1J6_3_LC_5_5_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 counter_RNIN1J6_3_LC_5_5_2 (
            .in0(_gnd_net_),
            .in1(N__20803),
            .in2(_gnd_net_),
            .in3(N__20791),
            .lcout(),
            .ltout(un2_counter_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIQKFG_5_LC_5_5_3.C_ON=1'b0;
    defparam counter_RNIQKFG_5_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam counter_RNIQKFG_5_LC_5_5_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNIQKFG_5_LC_5_5_3 (
            .in0(N__20779),
            .in1(N__20767),
            .in2(N__20756),
            .in3(N__20678),
            .lcout(un2_counter_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_12_LC_5_6_0.C_ON=1'b0;
    defparam counter_12_LC_5_6_0.SEQ_MODE=4'b1010;
    defparam counter_12_LC_5_6_0.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_12_LC_5_6_0 (
            .in0(N__21091),
            .in1(N__21058),
            .in2(N__20753),
            .in3(N__21023),
            .lcout(counterZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47999),
            .ce(),
            .sr(N__47329));
    defparam counter_10_LC_5_6_1.C_ON=1'b0;
    defparam counter_10_LC_5_6_1.SEQ_MODE=4'b1010;
    defparam counter_10_LC_5_6_1.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_10_LC_5_6_1 (
            .in0(N__21022),
            .in1(N__21090),
            .in2(N__20729),
            .in3(N__21059),
            .lcout(counterZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47999),
            .ce(),
            .sr(N__47329));
    defparam counter_1_LC_5_6_2.C_ON=1'b0;
    defparam counter_1_LC_5_6_2.SEQ_MODE=4'b1010;
    defparam counter_1_LC_5_6_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 counter_1_LC_5_6_2 (
            .in0(N__20685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20705),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47999),
            .ce(),
            .sr(N__47329));
    defparam counter_0_LC_5_6_4.C_ON=1'b0;
    defparam counter_0_LC_5_6_4.SEQ_MODE=4'b1010;
    defparam counter_0_LC_5_6_4.LUT_INIT=16'b0000011100001111;
    LogicCell40 counter_0_LC_5_6_4 (
            .in0(N__21089),
            .in1(N__21057),
            .in2(N__20687),
            .in3(N__21021),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47999),
            .ce(),
            .sr(N__47329));
    defparam \pwm_generator_inst.threshold_3_LC_5_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_5_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_5_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20660),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47998),
            .ce(),
            .sr(N__47342));
    defparam clk_10khz_LC_5_7_7.C_ON=1'b0;
    defparam clk_10khz_LC_5_7_7.SEQ_MODE=4'b1010;
    defparam clk_10khz_LC_5_7_7.LUT_INIT=16'b0111100011110000;
    LogicCell40 clk_10khz_LC_5_7_7 (
            .in0(N__21085),
            .in1(N__21055),
            .in2(N__22096),
            .in3(N__21025),
            .lcout(clk_10khz_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47998),
            .ce(),
            .sr(N__47342));
    defparam clk_10khz_RNIIENA2_LC_5_8_0.C_ON=1'b0;
    defparam clk_10khz_RNIIENA2_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam clk_10khz_RNIIENA2_LC_5_8_0.LUT_INIT=16'b0111100011110000;
    LogicCell40 clk_10khz_RNIIENA2_LC_5_8_0 (
            .in0(N__21084),
            .in1(N__21054),
            .in2(N__22092),
            .in3(N__21024),
            .lcout(clk_10khz_RNIIENAZ0Z2),
            .ltout(clk_10khz_RNIIENAZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_8_1 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__33693),
            .in2(N__20993),
            .in3(N__22085),
            .lcout(N_605_g),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_5_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_5_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_5_8_2  (
            .in0(N__20884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20845),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__27991),
            .in2(N__20978),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__27929),
            .in2(N__21947),
            .in3(N__20933),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__22001),
            .in2(N__30040),
            .in3(N__20915),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__27809),
            .in2(N__20912),
            .in3(N__20873),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__27754),
            .in2(N__21977),
            .in3(N__20834),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__27692),
            .in2(N__21359),
            .in3(N__21326),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__28517),
            .in2(N__25349),
            .in3(N__21296),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__21293),
            .in2(N__28448),
            .in3(N__21260),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__47992),
            .ce(N__32484),
            .sr(N__47360));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__28373),
            .in2(N__21257),
            .in3(N__21212),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__28303),
            .in2(N__25334),
            .in3(N__21173),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__28220),
            .in2(N__21170),
            .in3(N__21149),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__28145),
            .in2(N__21146),
            .in3(N__21122),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__28070),
            .in2(N__21119),
            .in3(N__21095),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__29056),
            .in2(N__21989),
            .in3(N__21518),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__28985),
            .in2(N__21959),
            .in3(N__21503),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__21500),
            .in2(N__28910),
            .in3(N__21482),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__47988),
            .ce(N__32432),
            .sr(N__47370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__21479),
            .in2(N__28841),
            .in3(N__21452),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__28751),
            .in2(N__22166),
            .in3(N__21437),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__28670),
            .in2(N__21434),
            .in3(N__21410),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__28592),
            .in2(N__21791),
            .in3(N__21395),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__29423),
            .in2(N__21392),
            .in3(N__21362),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__21725),
            .in2(N__29366),
            .in3(N__21704),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__29296),
            .in2(N__22181),
            .in3(N__21686),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__29222),
            .in2(N__22115),
            .in3(N__21674),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__47979),
            .ce(N__32489),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__21671),
            .in2(N__30407),
            .in3(N__21647),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__30356),
            .in2(N__22149),
            .in3(N__21629),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__22139),
            .in2(N__29114),
            .in3(N__21599),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__32596),
            .in2(N__22150),
            .in3(N__21578),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__22143),
            .in2(N__29705),
            .in3(N__21560),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__29636),
            .in2(N__22151),
            .in3(N__21542),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__22147),
            .in2(N__29576),
            .in3(N__21902),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7  (
            .in0(N__22148),
            .in1(N__33083),
            .in2(_gnd_net_),
            .in3(N__21899),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47969),
            .ce(N__32480),
            .sr(N__47382));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28555),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47961),
            .ce(N__32491),
            .sr(N__47390));
    defparam CONSTANT_ONE_LUT4_LC_5_28_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_28_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_28_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_6_LC_7_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_7_8_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_7_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21779),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_2_LC_7_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_7_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_7_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21770),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_0_LC_7_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_7_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21755),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_5_LC_7_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_7_8_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_7_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21746),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_7_LC_7_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_7_8_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_7_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21737),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_1_LC_7_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_7_8_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_7_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22049),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_4_LC_7_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_7_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_7_8_7  (
            .in0(N__22040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47989),
            .ce(),
            .sr(N__47330));
    defparam \pwm_generator_inst.threshold_9_LC_7_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22031),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47980),
            .ce(),
            .sr(N__47343));
    defparam \pwm_generator_inst.threshold_8_LC_7_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_7_9_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_7_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22016),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47980),
            .ce(),
            .sr(N__47343));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27859),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47970),
            .ce(N__32513),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29023),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47970),
            .ce(N__32513),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27721),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47970),
            .ce(N__32513),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28951),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47970),
            .ce(N__32513),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_7_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_7_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27895),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47970),
            .ce(N__32513),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_11_3  (
            .in0(N__29417),
            .in1(N__28591),
            .in2(N__29297),
            .in3(N__28747),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__27690),
            .in2(_gnd_net_),
            .in3(N__28441),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_7_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_7_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29257),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47956),
            .ce(N__32514),
            .sr(N__47371));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_7_12_1  (
            .in0(N__28708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47956),
            .ce(N__32514),
            .sr(N__47371));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29510),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47956),
            .ce(N__32514),
            .sr(N__47371));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29185),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47956),
            .ce(N__32514),
            .sr(N__47371));
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_13_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \current_shift_inst.phase_valid_RNISLOR2_LC_7_13_1  (
            .in0(N__30203),
            .in1(N__22100),
            .in2(N__33722),
            .in3(N__22064),
            .lcout(\current_shift_inst.phase_valid_RNISLORZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_21_LC_7_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_21_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_21_LC_7_14_5 .LUT_INIT=16'b1110110011111100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_21_LC_7_14_5  (
            .in0(N__22193),
            .in1(N__44200),
            .in2(N__39353),
            .in3(N__43963),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto31_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_7_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_7_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_7_15_0  (
            .in0(N__26489),
            .in1(N__27133),
            .in2(_gnd_net_),
            .in3(N__24913),
            .lcout(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_7_16_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__31231),
            .in2(_gnd_net_),
            .in3(N__31140),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_7_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_7_16_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__30596),
            .in2(_gnd_net_),
            .in3(N__30562),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_7_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_7_16_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_7_16_2  (
            .in0(N__31366),
            .in1(N__31141),
            .in2(N__31235),
            .in3(N__31336),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__30696),
            .in2(_gnd_net_),
            .in3(N__30656),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_4  (
            .in0(N__27043),
            .in1(N__23122),
            .in2(N__27011),
            .in3(N__27169),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__27042),
            .in2(_gnd_net_),
            .in3(N__27007),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_7_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_7_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_7_16_6  (
            .in0(N__30597),
            .in1(N__31271),
            .in2(N__30566),
            .in3(N__31189),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7  (
            .in0(N__27170),
            .in1(_gnd_net_),
            .in2(N__23126),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_7_17_0 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_7_17_0  (
            .in0(N__30845),
            .in1(N__25681),
            .in2(N__26648),
            .in3(N__30762),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_7_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_7_17_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_7_17_1  (
            .in0(N__25680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26643),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_7_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_7_17_2 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_7_17_2  (
            .in0(N__22639),
            .in1(N__27119),
            .in2(N__26456),
            .in3(N__24909),
            .lcout(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_7_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23339),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47919),
            .ce(N__22388),
            .sr(N__47398));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8SSQ5_15_LC_7_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8SSQ5_15_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8SSQ5_15_LC_7_17_4 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8SSQ5_15_LC_7_17_4  (
            .in0(N__42026),
            .in1(N__44156),
            .in2(N__42380),
            .in3(N__36845),
            .lcout(\delay_measurement_inst.delay_hc_reg3lt19_0 ),
            .ltout(\delay_measurement_inst.delay_hc_reg3lt19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_31_LC_7_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_31_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_31_LC_7_17_5 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_31_LC_7_17_5  (
            .in0(N__39352),
            .in1(N__44204),
            .in2(N__22184),
            .in3(N__43967),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_7_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_7_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_7_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23366),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47919),
            .ce(N__22388),
            .sr(N__47398));
    defparam \current_shift_inst.control_input_RNO_0_25_LC_7_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_7_18_2 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \current_shift_inst.control_input_RNO_0_25_LC_7_18_2  (
            .in0(N__27065),
            .in1(N__25297),
            .in2(N__27132),
            .in3(N__22741),
            .lcout(\current_shift_inst.un38_control_input_0_axb_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_18_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_18_3  (
            .in0(N__25027),
            .in1(N__22740),
            .in2(_gnd_net_),
            .in3(N__27064),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_7_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_7_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31931),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47913),
            .ce(N__31953),
            .sr(N__47402));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_7_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_7_18_6 .LUT_INIT=16'b0101010101100101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_7_18_6  (
            .in0(N__22611),
            .in1(N__22635),
            .in2(N__27131),
            .in3(N__24907),
            .lcout(\current_shift_inst.N_1620_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_7_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_7_18_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_7_18_7  (
            .in0(N__24908),
            .in1(N__22612),
            .in2(N__22640),
            .in3(N__27112),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_7_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_7_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_7_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__23362),
            .in2(N__23312),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_3 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_7_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__23335),
            .in2(N__23281),
            .in3(N__22217),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_7_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__23311),
            .in2(N__23254),
            .in3(N__22214),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_7_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__23224),
            .in2(N__23282),
            .in3(N__22211),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_7_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__23200),
            .in2(N__23255),
            .in3(N__22208),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_7_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__23225),
            .in2(N__23177),
            .in3(N__22205),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_7_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__23201),
            .in2(N__23612),
            .in3(N__22202),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_7_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_7_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__23176),
            .in2(N__23576),
            .in3(N__22199),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47907),
            .ce(N__22387),
            .sr(N__47405));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_7_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__23548),
            .in2(N__23611),
            .in3(N__22196),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_11 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_7_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__23575),
            .in2(N__23527),
            .in3(N__22244),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_7_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_7_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__23549),
            .in2(N__23500),
            .in3(N__22241),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_7_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_7_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__23467),
            .in2(N__23528),
            .in3(N__22238),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_7_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_7_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__23440),
            .in2(N__23501),
            .in3(N__22235),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_7_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_7_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__23416),
            .in2(N__23471),
            .in3(N__22232),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_7_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_7_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__23441),
            .in2(N__23396),
            .in3(N__22229),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_7_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_7_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__23417),
            .in2(N__23837),
            .in3(N__22226),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47902),
            .ce(N__22386),
            .sr(N__47408));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_7_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__23392),
            .in2(N__23804),
            .in3(N__22223),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_19 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_7_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__23770),
            .in2(N__23836),
            .in3(N__22220),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_7_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__23800),
            .in2(N__23746),
            .in3(N__22271),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_7_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__23771),
            .in2(N__23716),
            .in3(N__22268),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_7_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(N__23686),
            .in2(N__23747),
            .in3(N__22265),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_7_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__23662),
            .in2(N__23717),
            .in3(N__22262),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_7_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__23687),
            .in2(N__23642),
            .in3(N__22259),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_7_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_7_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_7_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__23663),
            .in2(N__24149),
            .in3(N__22256),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47895),
            .ce(N__22385),
            .sr(N__47412));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_7_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_7_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__23638),
            .in2(N__24113),
            .in3(N__22253),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_27 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47889),
            .ce(N__22384),
            .sr(N__47414));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_7_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_7_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_7_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(N__24082),
            .in2(N__24148),
            .in3(N__22250),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47889),
            .ce(N__22384),
            .sr(N__47414));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_7_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_7_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(N__24112),
            .in2(N__24062),
            .in3(N__22247),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47889),
            .ce(N__22384),
            .sr(N__47414));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_7_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_7_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__24083),
            .in2(N__24038),
            .in3(N__22394),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47889),
            .ce(N__22384),
            .sr(N__47414));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_7_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_7_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_7_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22391),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47889),
            .ce(N__22384),
            .sr(N__47414));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__22367),
            .in2(N__22361),
            .in3(N__24468),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__22352),
            .in2(N__22346),
            .in3(N__24384),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__22328),
            .in2(N__22337),
            .in3(N__24489),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__22307),
            .in2(N__22322),
            .in3(N__24405),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__22301),
            .in2(N__22295),
            .in3(N__24360),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__22286),
            .in2(N__22280),
            .in3(N__24315),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__22481),
            .in2(N__22475),
            .in3(N__24339),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__22457),
            .in2(N__22466),
            .in3(N__24213),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__22442),
            .in2(N__22451),
            .in3(N__24235),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__22427),
            .in2(N__22436),
            .in3(N__24255),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_8_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_8_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22421),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47971),
            .ce(),
            .sr(N__47331));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_0  (
            .in0(N__30041),
            .in1(N__27922),
            .in2(_gnd_net_),
            .in3(N__27992),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_8_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_8_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_8_10_1  (
            .in0(N__28984),
            .in1(N__28833),
            .in2(N__29057),
            .in3(N__28144),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_8_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_8_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_8_10_2  (
            .in0(N__29216),
            .in1(N__28906),
            .in2(N__29631),
            .in3(N__28212),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_8_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_8_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_8_10_4  (
            .in0(N__29694),
            .in1(N__32588),
            .in2(N__28069),
            .in3(N__29561),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA31P2_10_LC_8_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA31P2_10_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA31P2_10_LC_8_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA31P2_10_LC_8_10_5  (
            .in0(N__22535),
            .in1(N__22529),
            .in2(N__22523),
            .in3(N__22520),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_11_1  (
            .in0(N__28365),
            .in1(N__28509),
            .in2(N__28296),
            .in3(N__28440),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_11_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_11_2  (
            .in0(N__27760),
            .in1(N__27804),
            .in2(N__22514),
            .in3(N__27691),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_8_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_8_11_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_8_11_6  (
            .in0(N__28510),
            .in1(N__28366),
            .in2(N__28304),
            .in3(N__22511),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_8_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_8_11_7 .LUT_INIT=16'b1111001011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_8_11_7  (
            .in0(N__22505),
            .in1(N__27761),
            .in2(N__22499),
            .in3(N__27805),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_8_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_8_12_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_8_12_1  (
            .in0(N__36819),
            .in1(N__40724),
            .in2(_gnd_net_),
            .in3(N__22496),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47953),
            .ce(),
            .sr(N__47361));
    defparam \current_shift_inst.control_input_0_LC_8_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__24608),
            .in2(N__29948),
            .in3(N__29947),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_8_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__24599),
            .in2(_gnd_net_),
            .in3(N__22487),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_8_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_8_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__24590),
            .in2(_gnd_net_),
            .in3(N__22484),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_8_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__24581),
            .in2(_gnd_net_),
            .in3(N__22562),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_8_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_8_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__24572),
            .in2(_gnd_net_),
            .in3(N__22559),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_8_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_8_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__24563),
            .in2(_gnd_net_),
            .in3(N__22556),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_8_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_8_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__24713),
            .in2(_gnd_net_),
            .in3(N__22553),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_8_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__24692),
            .in2(_gnd_net_),
            .in3(N__22550),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__47944),
            .ce(N__24952),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_8_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_8_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__24671),
            .in2(_gnd_net_),
            .in3(N__22547),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_8_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_8_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__24662),
            .in2(_gnd_net_),
            .in3(N__22544),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_8_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_8_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__24653),
            .in2(_gnd_net_),
            .in3(N__22541),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_8_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_11_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_8_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_11_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__24644),
            .in2(_gnd_net_),
            .in3(N__22538),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_10 ),
            .carryout(\current_shift_inst.control_input_1_cry_11 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_12_LC_8_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_12_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_12_LC_8_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_12_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__24635),
            .in2(_gnd_net_),
            .in3(N__22589),
            .lcout(\current_shift_inst.control_inputZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_11 ),
            .carryout(\current_shift_inst.control_input_1_cry_12 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_13_LC_8_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_13_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_13_LC_8_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_13_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__24626),
            .in2(_gnd_net_),
            .in3(N__22586),
            .lcout(\current_shift_inst.control_inputZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_12 ),
            .carryout(\current_shift_inst.control_input_1_cry_13 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_14_LC_8_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_14_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_14_LC_8_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_14_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__24617),
            .in2(_gnd_net_),
            .in3(N__22583),
            .lcout(\current_shift_inst.control_inputZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_13 ),
            .carryout(\current_shift_inst.control_input_1_cry_14 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_15_LC_8_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_15_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_15_LC_8_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_15_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__24839),
            .in2(_gnd_net_),
            .in3(N__22580),
            .lcout(\current_shift_inst.control_inputZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_14 ),
            .carryout(\current_shift_inst.control_input_1_cry_15 ),
            .clk(N__47935),
            .ce(N__24968),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_16_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_16_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_16_LC_8_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_16_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__24830),
            .in2(_gnd_net_),
            .in3(N__22577),
            .lcout(\current_shift_inst.control_inputZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.control_input_1_cry_16 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_17_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_17_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_17_LC_8_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_17_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__24821),
            .in2(_gnd_net_),
            .in3(N__22574),
            .lcout(\current_shift_inst.control_inputZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_16 ),
            .carryout(\current_shift_inst.control_input_1_cry_17 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_18_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_18_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_18_LC_8_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_18_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__24791),
            .in2(_gnd_net_),
            .in3(N__22571),
            .lcout(\current_shift_inst.control_inputZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_17 ),
            .carryout(\current_shift_inst.control_input_1_cry_18 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_19_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_19_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_19_LC_8_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_19_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__24782),
            .in2(_gnd_net_),
            .in3(N__22568),
            .lcout(\current_shift_inst.control_inputZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_18 ),
            .carryout(\current_shift_inst.control_input_1_cry_19 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_20_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_20_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_20_LC_8_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_20_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__24752),
            .in2(_gnd_net_),
            .in3(N__22565),
            .lcout(\current_shift_inst.control_inputZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_19 ),
            .carryout(\current_shift_inst.control_input_1_cry_20 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_21_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_21_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_21_LC_8_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_21_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__24743),
            .in2(_gnd_net_),
            .in3(N__22655),
            .lcout(\current_shift_inst.control_inputZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_20 ),
            .carryout(\current_shift_inst.control_input_1_cry_21 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_22_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_22_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_22_LC_8_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_22_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__24722),
            .in2(_gnd_net_),
            .in3(N__22652),
            .lcout(\current_shift_inst.control_inputZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_21 ),
            .carryout(\current_shift_inst.control_input_1_cry_22 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_23_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_23_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_23_LC_8_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_23_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__25049),
            .in2(_gnd_net_),
            .in3(N__22649),
            .lcout(\current_shift_inst.control_inputZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_22 ),
            .carryout(\current_shift_inst.control_input_1_cry_23 ),
            .clk(N__47926),
            .ce(N__24959),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_24_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_24_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_24_LC_8_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_24_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__25001),
            .in2(_gnd_net_),
            .in3(N__22646),
            .lcout(\current_shift_inst.control_inputZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_24 ),
            .clk(N__47920),
            .ce(N__24966),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22643),
            .lcout(\current_shift_inst.control_input_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__24900),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.z_5_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_8_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__22634),
            .in2(N__23032),
            .in3(N__22616),
            .lcout(\current_shift_inst.z_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_1 ),
            .carryout(\current_shift_inst.z_5_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_8_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__22613),
            .in2(N__23035),
            .in3(N__22595),
            .lcout(\current_shift_inst.z_5_3 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_2 ),
            .carryout(\current_shift_inst.z_5_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_8_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__25590),
            .in2(N__23033),
            .in3(N__22592),
            .lcout(\current_shift_inst.z_5_4 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_3 ),
            .carryout(\current_shift_inst.z_5_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__25630),
            .in2(N__23036),
            .in3(N__22682),
            .lcout(\current_shift_inst.z_5_5 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_4 ),
            .carryout(\current_shift_inst.z_5_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__25488),
            .in2(N__23034),
            .in3(N__22679),
            .lcout(\current_shift_inst.z_5_6 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_5 ),
            .carryout(\current_shift_inst.z_5_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__22967),
            .in2(N__25880),
            .in3(N__22676),
            .lcout(\current_shift_inst.z_5_7 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_6 ),
            .carryout(\current_shift_inst.z_5_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__22974),
            .in2(N__25739),
            .in3(N__22673),
            .lcout(\current_shift_inst.z_5_8 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_7 ),
            .carryout(\current_shift_inst.z_5_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_8_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__25753),
            .in2(N__23088),
            .in3(N__22670),
            .lcout(\current_shift_inst.z_5_9 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.z_5_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_8_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__25909),
            .in2(N__23084),
            .in3(N__22667),
            .lcout(\current_shift_inst.z_5_10 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_9 ),
            .carryout(\current_shift_inst.z_5_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_8_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__30867),
            .in2(N__23086),
            .in3(N__22664),
            .lcout(\current_shift_inst.z_5_11 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_10 ),
            .carryout(\current_shift_inst.z_5_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_8_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__30746),
            .in2(N__23085),
            .in3(N__22661),
            .lcout(\current_shift_inst.z_5_12 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_11 ),
            .carryout(\current_shift_inst.z_5_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_8_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__25676),
            .in2(N__23087),
            .in3(N__22658),
            .lcout(\current_shift_inst.z_5_13 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_12 ),
            .carryout(\current_shift_inst.z_5_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_8_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__23050),
            .in2(N__25826),
            .in3(N__22709),
            .lcout(\current_shift_inst.z_5_14 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_13 ),
            .carryout(\current_shift_inst.z_5_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_8_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__23043),
            .in2(N__26139),
            .in3(N__22706),
            .lcout(\current_shift_inst.z_5_15 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_14 ),
            .carryout(\current_shift_inst.z_5_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_8_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_8_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__23051),
            .in2(N__26187),
            .in3(N__22703),
            .lcout(\current_shift_inst.z_5_16 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_15 ),
            .carryout(\current_shift_inst.z_5_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_8_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__26005),
            .in2(N__23027),
            .in3(N__22700),
            .lcout(\current_shift_inst.z_5_17 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.z_5_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_8_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__25971),
            .in2(N__23030),
            .in3(N__22697),
            .lcout(\current_shift_inst.z_5_18 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_17 ),
            .carryout(\current_shift_inst.z_5_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_8_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__26218),
            .in2(N__23028),
            .in3(N__22694),
            .lcout(\current_shift_inst.z_5_19 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_18 ),
            .carryout(\current_shift_inst.z_5_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_8_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__26086),
            .in2(N__23031),
            .in3(N__22691),
            .lcout(\current_shift_inst.z_5_20 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_19 ),
            .carryout(\current_shift_inst.z_5_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_8_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__26049),
            .in2(N__23029),
            .in3(N__22688),
            .lcout(\current_shift_inst.z_5_21 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_20 ),
            .carryout(\current_shift_inst.z_5_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_8_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__22949),
            .in2(N__30506),
            .in3(N__22685),
            .lcout(\current_shift_inst.z_5_22 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_21 ),
            .carryout(\current_shift_inst.z_5_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__22957),
            .in2(N__30598),
            .in3(N__23144),
            .lcout(\current_shift_inst.z_5_23 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_22 ),
            .carryout(\current_shift_inst.z_5_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__22950),
            .in2(N__31275),
            .in3(N__23141),
            .lcout(\current_shift_inst.z_5_24 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_23 ),
            .carryout(\current_shift_inst.z_5_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_8_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__31128),
            .in2(N__22874),
            .in3(N__23138),
            .lcout(\current_shift_inst.z_5_25 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.z_5_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__31353),
            .in2(N__22877),
            .in3(N__23135),
            .lcout(\current_shift_inst.z_5_26 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_25 ),
            .carryout(\current_shift_inst.z_5_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__30683),
            .in2(N__22875),
            .in3(N__23132),
            .lcout(\current_shift_inst.z_5_27 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_26 ),
            .carryout(\current_shift_inst.z_5_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__27038),
            .in2(N__22878),
            .in3(N__23129),
            .lcout(\current_shift_inst.z_5_28 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_27 ),
            .carryout(\current_shift_inst.z_5_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_8_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__23121),
            .in2(N__22876),
            .in3(N__23102),
            .lcout(\current_shift_inst.z_5_29 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_28 ),
            .carryout(\current_shift_inst.z_5_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_8_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__22838),
            .in2(N__22742),
            .in3(N__22715),
            .lcout(\current_shift_inst.z_5_30 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_29 ),
            .carryout(\current_shift_inst.z_5_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_8_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_8_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22712),
            .lcout(\current_shift_inst.z_5_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.counter_0_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_0_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_0_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_0_LC_8_21_0  (
            .in0(N__23955),
            .in1(N__23355),
            .in2(_gnd_net_),
            .in3(N__23342),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_0 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_1_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_1_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_1_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_1_LC_8_21_1  (
            .in0(N__23950),
            .in1(N__23328),
            .in2(_gnd_net_),
            .in3(N__23315),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_1 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_2_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_2_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_2_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_2_LC_8_21_2  (
            .in0(N__23956),
            .in1(N__23307),
            .in2(_gnd_net_),
            .in3(N__23285),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_2 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_3_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_3_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_3_LC_8_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_3_LC_8_21_3  (
            .in0(N__23951),
            .in1(N__23274),
            .in2(_gnd_net_),
            .in3(N__23258),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_3 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_4_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_4_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_4_LC_8_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_4_LC_8_21_4  (
            .in0(N__23957),
            .in1(N__23242),
            .in2(_gnd_net_),
            .in3(N__23228),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_4 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_5_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_5_LC_8_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_5_LC_8_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_5_LC_8_21_5  (
            .in0(N__23952),
            .in1(N__23218),
            .in2(_gnd_net_),
            .in3(N__23204),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_5 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_6_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_6_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_6_LC_8_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_6_LC_8_21_6  (
            .in0(N__23954),
            .in1(N__23194),
            .in2(_gnd_net_),
            .in3(N__23180),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_6 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_7_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_7_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_7_LC_8_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_7_LC_8_21_7  (
            .in0(N__23953),
            .in1(N__23161),
            .in2(_gnd_net_),
            .in3(N__23147),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_7 ),
            .clk(N__47890),
            .ce(N__24005),
            .sr(N__47409));
    defparam \current_shift_inst.timer_phase.counter_8_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_8_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_8_LC_8_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_8_LC_8_22_0  (
            .in0(N__23949),
            .in1(N__23601),
            .in2(_gnd_net_),
            .in3(N__23579),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_8 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_9_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_9_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_9_LC_8_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_9_LC_8_22_1  (
            .in0(N__23961),
            .in1(N__23571),
            .in2(_gnd_net_),
            .in3(N__23552),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_9 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_10_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_10_LC_8_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_10_LC_8_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_10_LC_8_22_2  (
            .in0(N__23946),
            .in1(N__23547),
            .in2(_gnd_net_),
            .in3(N__23531),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_10 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_11_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_11_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_11_LC_8_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_11_LC_8_22_3  (
            .in0(N__23958),
            .in1(N__23520),
            .in2(_gnd_net_),
            .in3(N__23504),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_11 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_12_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_12_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_12_LC_8_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_12_LC_8_22_4  (
            .in0(N__23947),
            .in1(N__23488),
            .in2(_gnd_net_),
            .in3(N__23474),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_12 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_13_LC_8_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_13_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_13_LC_8_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_13_LC_8_22_5  (
            .in0(N__23959),
            .in1(N__23460),
            .in2(_gnd_net_),
            .in3(N__23444),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_13 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_14_LC_8_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_14_LC_8_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_14_LC_8_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_14_LC_8_22_6  (
            .in0(N__23948),
            .in1(N__23434),
            .in2(_gnd_net_),
            .in3(N__23420),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_14 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_15_LC_8_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_15_LC_8_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_15_LC_8_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_15_LC_8_22_7  (
            .in0(N__23960),
            .in1(N__23415),
            .in2(_gnd_net_),
            .in3(N__23399),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_15 ),
            .clk(N__47884),
            .ce(N__24000),
            .sr(N__47413));
    defparam \current_shift_inst.timer_phase.counter_16_LC_8_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_16_LC_8_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_16_LC_8_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_16_LC_8_23_0  (
            .in0(N__23962),
            .in1(N__23388),
            .in2(_gnd_net_),
            .in3(N__23369),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_23_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_16 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_17_LC_8_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_17_LC_8_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_17_LC_8_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_17_LC_8_23_1  (
            .in0(N__23966),
            .in1(N__23826),
            .in2(_gnd_net_),
            .in3(N__23807),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_17 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_18_LC_8_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_18_LC_8_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_18_LC_8_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_18_LC_8_23_2  (
            .in0(N__23963),
            .in1(N__23799),
            .in2(_gnd_net_),
            .in3(N__23774),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_18 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_19_LC_8_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_19_LC_8_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_19_LC_8_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_19_LC_8_23_3  (
            .in0(N__23967),
            .in1(N__23769),
            .in2(_gnd_net_),
            .in3(N__23750),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_19 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_20_LC_8_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_20_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_20_LC_8_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_20_LC_8_23_4  (
            .in0(N__23964),
            .in1(N__23734),
            .in2(_gnd_net_),
            .in3(N__23720),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_20 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_21_LC_8_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_21_LC_8_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_21_LC_8_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_21_LC_8_23_5  (
            .in0(N__23968),
            .in1(N__23704),
            .in2(_gnd_net_),
            .in3(N__23690),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_21 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_22_LC_8_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_22_LC_8_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_22_LC_8_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_22_LC_8_23_6  (
            .in0(N__23965),
            .in1(N__23680),
            .in2(_gnd_net_),
            .in3(N__23666),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_22 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_23_LC_8_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_23_LC_8_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_23_LC_8_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_23_LC_8_23_7  (
            .in0(N__23969),
            .in1(N__23661),
            .in2(_gnd_net_),
            .in3(N__23645),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_23 ),
            .clk(N__47881),
            .ce(N__24001),
            .sr(N__47415));
    defparam \current_shift_inst.timer_phase.counter_24_LC_8_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_24_LC_8_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_24_LC_8_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_24_LC_8_24_0  (
            .in0(N__23940),
            .in1(N__23634),
            .in2(_gnd_net_),
            .in3(N__23615),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_24_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_24 ),
            .clk(N__47875),
            .ce(N__23985),
            .sr(N__47417));
    defparam \current_shift_inst.timer_phase.counter_25_LC_8_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_25_LC_8_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_25_LC_8_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_25_LC_8_24_1  (
            .in0(N__23944),
            .in1(N__24135),
            .in2(_gnd_net_),
            .in3(N__24116),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_25 ),
            .clk(N__47875),
            .ce(N__23985),
            .sr(N__47417));
    defparam \current_shift_inst.timer_phase.counter_26_LC_8_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_26_LC_8_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_26_LC_8_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_26_LC_8_24_2  (
            .in0(N__23941),
            .in1(N__24108),
            .in2(_gnd_net_),
            .in3(N__24086),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_26 ),
            .clk(N__47875),
            .ce(N__23985),
            .sr(N__47417));
    defparam \current_shift_inst.timer_phase.counter_27_LC_8_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_27_LC_8_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_27_LC_8_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_27_LC_8_24_3  (
            .in0(N__23945),
            .in1(N__24081),
            .in2(_gnd_net_),
            .in3(N__24065),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_27 ),
            .clk(N__47875),
            .ce(N__23985),
            .sr(N__47417));
    defparam \current_shift_inst.timer_phase.counter_28_LC_8_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_28_LC_8_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_28_LC_8_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_28_LC_8_24_4  (
            .in0(N__23942),
            .in1(N__24058),
            .in2(_gnd_net_),
            .in3(N__24044),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_28 ),
            .clk(N__47875),
            .ce(N__23985),
            .sr(N__47417));
    defparam \current_shift_inst.timer_phase.counter_29_LC_8_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.counter_29_LC_8_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_29_LC_8_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_phase.counter_29_LC_8_24_5  (
            .in0(N__24034),
            .in1(N__23943),
            .in2(_gnd_net_),
            .in3(N__24041),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47875),
            .ce(N__23985),
            .sr(N__47417));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_8_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_8_25_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_8_25_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_8_25_1  (
            .in0(_gnd_net_),
            .in1(N__27563),
            .in2(_gnd_net_),
            .in3(N__27539),
            .lcout(\current_shift_inst.timer_s1.N_187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_8_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_8_25_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_8_25_2 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIL91O_LC_8_25_2  (
            .in0(N__27472),
            .in1(N__25263),
            .in2(_gnd_net_),
            .in3(N__27452),
            .lcout(\current_shift_inst.timer_phase.N_193_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_8_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_8_25_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_8_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIB31B_LC_8_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27471),
            .lcout(\current_shift_inst.timer_phase.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_4_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_4_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_9_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23849),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47995),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_9_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_9_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_9_7_0  (
            .in0(N__24296),
            .in1(N__24469),
            .in2(_gnd_net_),
            .in3(N__24176),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_1_LC_9_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_9_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_9_7_1  (
            .in0(N__24292),
            .in1(N__24388),
            .in2(_gnd_net_),
            .in3(N__24173),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_2_LC_9_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_9_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_9_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_9_7_2  (
            .in0(N__24297),
            .in1(N__24490),
            .in2(_gnd_net_),
            .in3(N__24170),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_3_LC_9_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_9_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_9_7_3  (
            .in0(N__24293),
            .in1(N__24409),
            .in2(_gnd_net_),
            .in3(N__24167),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_4_LC_9_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_9_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_9_7_4  (
            .in0(N__24298),
            .in1(N__24364),
            .in2(_gnd_net_),
            .in3(N__24164),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_5_LC_9_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_9_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_9_7_5  (
            .in0(N__24294),
            .in1(N__24316),
            .in2(_gnd_net_),
            .in3(N__24161),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_6_LC_9_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_9_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_9_7_6  (
            .in0(N__24299),
            .in1(N__24340),
            .in2(_gnd_net_),
            .in3(N__24158),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_7_LC_9_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_9_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_9_7_7  (
            .in0(N__24295),
            .in1(N__24217),
            .in2(_gnd_net_),
            .in3(N__24155),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__47981),
            .ce(),
            .sr(N__47310));
    defparam \pwm_generator_inst.counter_8_LC_9_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_9_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_9_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_9_8_0  (
            .in0(N__24291),
            .in1(N__24236),
            .in2(_gnd_net_),
            .in3(N__24152),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__47972),
            .ce(),
            .sr(N__47316));
    defparam \pwm_generator_inst.counter_9_LC_9_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_9_8_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_9_8_1  (
            .in0(N__24256),
            .in1(N__24290),
            .in2(_gnd_net_),
            .in3(N__24413),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47972),
            .ce(),
            .sr(N__47316));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_9_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_9_9_1 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_9_9_1  (
            .in0(N__24410),
            .in1(N__24389),
            .in2(N__24368),
            .in3(N__24449),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_9_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_9_9_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_9_9_2  (
            .in0(N__24197),
            .in1(N__24344),
            .in2(N__24323),
            .in3(N__24320),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_9_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_9_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_9_9_5  (
            .in0(N__24257),
            .in1(N__24234),
            .in2(_gnd_net_),
            .in3(N__24218),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3MVS6_31_LC_9_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3MVS6_31_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3MVS6_31_LC_9_9_7 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3MVS6_31_LC_9_9_7  (
            .in0(N__33069),
            .in1(N__30104),
            .in2(_gnd_net_),
            .in3(N__30075),
            .lcout(\current_shift_inst.PI_CTRL.N_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_9_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_9_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_9_10_0  (
            .in0(N__29615),
            .in1(N__28901),
            .in2(N__28219),
            .in3(N__29217),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI775B_18_LC_9_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI775B_18_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI775B_18_LC_9_10_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI775B_18_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__33011),
            .in2(_gnd_net_),
            .in3(N__28655),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_9_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_9_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_9_10_3  (
            .in0(N__29693),
            .in1(N__32589),
            .in2(N__29568),
            .in3(N__28056),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI50UD2_10_LC_9_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI50UD2_10_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI50UD2_10_LC_9_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI50UD2_10_LC_9_10_4  (
            .in0(N__24497),
            .in1(N__24191),
            .in2(N__24185),
            .in3(N__24182),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_9_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_9_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_9_10_6  (
            .in0(N__28979),
            .in1(N__29046),
            .in2(N__28837),
            .in3(N__28133),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_9_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_9_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_9_10_7  (
            .in0(N__24491),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24470),
            .lcout(\pwm_generator_inst.un1_counterlto2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_9_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_9_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_9_11_1  (
            .in0(N__30347),
            .in1(N__30392),
            .in2(N__29100),
            .in3(N__29354),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIO0BU3_18_LC_9_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIO0BU3_18_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIO0BU3_18_LC_9_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIO0BU3_18_LC_9_11_2  (
            .in0(N__33062),
            .in1(N__28659),
            .in2(N__24443),
            .in3(N__24440),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_9_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_9_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_9_11_4  (
            .in0(N__29355),
            .in1(N__30348),
            .in2(N__30402),
            .in3(N__29093),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_9_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_9_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_9_11_5  (
            .in0(N__29418),
            .in1(N__28736),
            .in2(N__29292),
            .in3(N__28583),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_17_LC_9_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_17_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_17_LC_9_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_17_LC_9_11_6  (
            .in0(N__24434),
            .in1(N__24428),
            .in2(N__24422),
            .in3(N__24419),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_12_0 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_9_12_0  (
            .in0(N__33063),
            .in1(N__32826),
            .in2(N__28688),
            .in3(N__32703),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47945),
            .ce(N__32549),
            .sr(N__47353));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_12_2 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_9_12_2  (
            .in0(N__33066),
            .in1(N__32835),
            .in2(N__29528),
            .in3(N__32708),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47945),
            .ce(N__32549),
            .sr(N__47353));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_4 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_4  (
            .in0(N__33064),
            .in1(N__32830),
            .in2(N__29384),
            .in3(N__32705),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47945),
            .ce(N__32549),
            .sr(N__47353));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5  (
            .in0(N__32706),
            .in1(N__29234),
            .in2(N__32864),
            .in3(N__33068),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47945),
            .ce(N__32549),
            .sr(N__47353));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6  (
            .in0(N__33065),
            .in1(N__32834),
            .in2(N__29162),
            .in3(N__32707),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47945),
            .ce(N__32549),
            .sr(N__47353));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_12_7 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_9_12_7  (
            .in0(N__32704),
            .in1(N__28529),
            .in2(N__32863),
            .in3(N__33067),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47945),
            .ce(N__32549),
            .sr(N__47353));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__27142),
            .in2(N__27146),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__24554),
            .in2(N__26510),
            .in3(N__29972),
            .lcout(\current_shift_inst.z_i_0_31 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__26488),
            .in2(N__24548),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__26455),
            .in2(N__24533),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_1 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4  (
            .in0(N__24518),
            .in1(N__26420),
            .in2(N__24506),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_2 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__25433),
            .in2(N__25459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_3 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__25568),
            .in2(N__25427),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_4 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__25415),
            .in2(N__25370),
            .in3(N__24602),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_5 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__25511),
            .in2(N__25469),
            .in3(N__24593),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__25847),
            .in2(N__25523),
            .in3(N__24584),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_7 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__25706),
            .in2(N__25397),
            .in3(N__24575),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_8 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__25898),
            .in2(N__25379),
            .in3(N__24566),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_9 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__25949),
            .in2(N__25550),
            .in3(N__24557),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_10 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__30725),
            .in2(N__25406),
            .in3(N__24707),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_11 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__24704),
            .in2(N__25388),
            .in3(N__24686),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_12 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__24683),
            .in2(N__25652),
            .in3(N__24665),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_13 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__25529),
            .in2(N__25793),
            .in3(N__24656),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__26108),
            .in2(N__25559),
            .in3(N__24647),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_15 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__26156),
            .in2(N__25538),
            .in3(N__24638),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_16 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__25955),
            .in2(N__26258),
            .in3(N__24629),
            .lcout(\current_shift_inst.control_input_1_axb_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_17 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__25700),
            .in2(N__26267),
            .in3(N__24620),
            .lcout(\current_shift_inst.control_input_1_axb_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_18 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__26201),
            .in2(N__25943),
            .in3(N__24611),
            .lcout(\current_shift_inst.control_input_1_axb_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_19 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__26030),
            .in2(N__26249),
            .in3(N__24833),
            .lcout(\current_shift_inst.control_input_1_axb_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_20 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__25694),
            .in2(N__26276),
            .in3(N__24824),
            .lcout(\current_shift_inst.control_input_1_axb_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_21 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__30527),
            .in2(N__30434),
            .in3(N__24815),
            .lcout(\current_shift_inst.control_input_1_axb_17 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__24812),
            .in2(N__24803),
            .in3(N__24785),
            .lcout(\current_shift_inst.control_input_1_axb_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_23 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__31112),
            .in2(N__30713),
            .in3(N__24776),
            .lcout(\current_shift_inst.control_input_1_axb_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_24 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__24773),
            .in2(N__24764),
            .in3(N__24746),
            .lcout(\current_shift_inst.control_input_1_axb_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_25 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__30614),
            .in2(N__31298),
            .in3(N__24737),
            .lcout(\current_shift_inst.control_input_1_axb_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_26 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__26978),
            .in2(N__24734),
            .in3(N__24716),
            .lcout(\current_shift_inst.control_input_1_axb_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_27 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__25070),
            .in2(N__25061),
            .in3(N__25043),
            .lcout(\current_shift_inst.control_input_1_axb_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_28 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__25040),
            .in2(N__25028),
            .in3(N__24995),
            .lcout(\current_shift_inst.control_input_1_axb_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_29 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_25_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_25_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_25_LC_9_17_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.control_input_25_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__24992),
            .in2(N__24980),
            .in3(N__24971),
            .lcout(\current_shift_inst.control_inputZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47908),
            .ce(N__24967),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_9_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__26500),
            .in2(N__24923),
            .in3(N__29768),
            .lcout(G_406),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.z_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_9_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__26475),
            .in2(N__24875),
            .in3(N__24914),
            .lcout(G_405),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_0 ),
            .carryout(\current_shift_inst.z_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_9_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_2_c_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__24866),
            .in2(N__26448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_1 ),
            .carryout(\current_shift_inst.z_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_9_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_3_c_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__26413),
            .in2(N__24857),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_2 ),
            .carryout(\current_shift_inst.z_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_9_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_4_c_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__26388),
            .in2(N__24848),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_3 ),
            .carryout(\current_shift_inst.z_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_9_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_5_c_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__25124),
            .in2(N__26366),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_4 ),
            .carryout(\current_shift_inst.z_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_9_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_6_c_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__25118),
            .in2(N__26336),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_5 ),
            .carryout(\current_shift_inst.z_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_9_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_7_c_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__25112),
            .in2(N__26303),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_6 ),
            .carryout(\current_shift_inst.z_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_8_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__25106),
            .in2(N__26765),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.z_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_9_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_9_c_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25097),
            .in2(N__26720),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_8 ),
            .carryout(\current_shift_inst.z_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_9_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_10_c_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__25091),
            .in2(N__26681),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_9 ),
            .carryout(\current_shift_inst.z_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_9_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_11_c_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__25085),
            .in2(N__30797),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_10 ),
            .carryout(\current_shift_inst.z_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_9_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_12_c_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__30827),
            .in2(N__25079),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_11 ),
            .carryout(\current_shift_inst.z_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_9_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_13_c_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__25184),
            .in2(N__26634),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_12 ),
            .carryout(\current_shift_inst.z_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_9_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_14_c_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__25178),
            .in2(N__26597),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_13 ),
            .carryout(\current_shift_inst.z_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_9_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_15_c_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__26556),
            .in2(N__25172),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_14 ),
            .carryout(\current_shift_inst.z_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_9_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_16_c_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__26524),
            .in2(N__25163),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.z_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_9_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_17_c_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__25148),
            .in2(N__26951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_16 ),
            .carryout(\current_shift_inst.z_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_9_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_18_c_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__25142),
            .in2(N__26912),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_17 ),
            .carryout(\current_shift_inst.z_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_9_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_19_c_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__25136),
            .in2(N__26868),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_18 ),
            .carryout(\current_shift_inst.z_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_9_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_20_c_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__25130),
            .in2(N__26840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_19 ),
            .carryout(\current_shift_inst.z_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_9_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_21_c_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__26799),
            .in2(N__25247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_20 ),
            .carryout(\current_shift_inst.z_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_9_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_22_c_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__25238),
            .in2(N__30459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_21 ),
            .carryout(\current_shift_inst.z_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_9_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_23_c_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__25232),
            .in2(N__30552),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_22 ),
            .carryout(\current_shift_inst.z_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_9_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_24_c_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__25226),
            .in2(N__31178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.z_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_9_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_25_c_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__25217),
            .in2(N__31220),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_24 ),
            .carryout(\current_shift_inst.z_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_9_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_26_c_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__25211),
            .in2(N__31323),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_25 ),
            .carryout(\current_shift_inst.z_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_9_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_27_c_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__25205),
            .in2(N__30644),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_26 ),
            .carryout(\current_shift_inst.z_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_9_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_28_c_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__25199),
            .in2(N__27001),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_27 ),
            .carryout(\current_shift_inst.z_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_9_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_29_c_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__27160),
            .in2(N__25193),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_28 ),
            .carryout(\current_shift_inst.z_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_9_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_9_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_30_c_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__27055),
            .in2(N__25316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_29 ),
            .carryout(\current_shift_inst.z_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_9_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_9_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.un10_control_input_z_s_31_LC_9_21_7  (
            .in0(N__27135),
            .in1(N__25307),
            .in2(N__25301),
            .in3(N__25277),
            .lcout(\current_shift_inst.z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_9_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_9_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.stop_timer_s1_RNO_0_LC_9_23_2  (
            .in0(N__30198),
            .in1(N__30278),
            .in2(N__27614),
            .in3(N__30245),
            .lcout(\current_shift_inst.stop_timer_s1_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_LC_9_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_9_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_9_24_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_9_24_1  (
            .in0(N__27602),
            .in1(N__27568),
            .in2(_gnd_net_),
            .in3(N__27541),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47868),
            .ce(),
            .sr(N__47416));
    defparam \current_shift_inst.meas_state_0_LC_9_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.meas_state_0_LC_9_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.meas_state_0_LC_9_24_3 .LUT_INIT=16'b0111111111001100;
    LogicCell40 \current_shift_inst.meas_state_0_LC_9_24_3  (
            .in0(N__30202),
            .in1(N__30279),
            .in2(N__27612),
            .in3(N__30244),
            .lcout(\current_shift_inst.meas_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47868),
            .ce(),
            .sr(N__47416));
    defparam \current_shift_inst.start_timer_phase_LC_9_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_phase_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_phase_LC_9_25_0 .LUT_INIT=16'b0011101100101010;
    LogicCell40 \current_shift_inst.start_timer_phase_LC_9_25_0  (
            .in0(N__25265),
            .in1(N__30281),
            .in2(N__32306),
            .in3(N__30246),
            .lcout(\current_shift_inst.start_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(N__35837),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_9_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_9_25_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_s1_LC_9_25_6 .LUT_INIT=16'b0111001111110000;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_9_25_6  (
            .in0(N__30194),
            .in1(N__30280),
            .in2(N__27613),
            .in3(N__30247),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(N__35837),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_9_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_s1_LC_9_25_7 .LUT_INIT=16'b1111110111001100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_9_25_7  (
            .in0(N__30248),
            .in1(N__25274),
            .in2(N__30289),
            .in3(N__27542),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(N__35837),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_LC_9_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_LC_9_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.running_LC_9_26_5 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_phase.running_LC_9_26_5  (
            .in0(N__25264),
            .in1(N__27473),
            .in2(_gnd_net_),
            .in3(N__27450),
            .lcout(\current_shift_inst.timer_phase.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47857),
            .ce(),
            .sr(N__47422));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_7_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_7_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25358),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47963),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28483),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47955),
            .ce(N__32550),
            .sr(N__47311));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_10_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_10_9_5 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_10_9_5  (
            .in0(N__33074),
            .in1(N__32881),
            .in2(N__28385),
            .in3(N__32638),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47955),
            .ce(N__32550),
            .sr(N__47311));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28265),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47955),
            .ce(N__32550),
            .sr(N__47311));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_10_0 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_10_10_0  (
            .in0(N__33036),
            .in1(N__32838),
            .in2(N__28607),
            .in3(N__32656),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_10_1 .LUT_INIT=16'b1111000111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_10_10_1  (
            .in0(N__30117),
            .in1(N__32842),
            .in2(N__27773),
            .in3(N__30074),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_10_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_10_10_2 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_10_10_2  (
            .in0(N__33034),
            .in1(N__32836),
            .in2(N__28997),
            .in3(N__32653),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_10_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_10_10_3 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_10_10_3  (
            .in0(N__32655),
            .in1(N__28850),
            .in2(N__33073),
            .in3(N__32839),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_10_4 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_10_10_4  (
            .in0(N__33035),
            .in1(N__32837),
            .in2(N__28925),
            .in3(N__32654),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_10_5 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_10_10_5  (
            .in0(N__30116),
            .in1(N__32840),
            .in2(N__27875),
            .in3(N__30073),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_10_7 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_10_10_7  (
            .in0(N__32657),
            .in1(N__33037),
            .in2(N__29594),
            .in3(N__32841),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47946),
            .ce(N__32553),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_11_0 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_10_11_0  (
            .in0(N__32714),
            .in1(N__28457),
            .in2(N__32861),
            .in3(N__33081),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_11_1 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_10_11_1  (
            .in0(N__33076),
            .in1(N__32811),
            .in2(N__28082),
            .in3(N__32710),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_11_2 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_10_11_2  (
            .in0(N__32711),
            .in1(N__28004),
            .in2(N__32859),
            .in3(N__33079),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_11_3 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_10_11_3  (
            .in0(N__33078),
            .in1(N__32825),
            .in2(N__28232),
            .in3(N__32716),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_11_4 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_10_11_4  (
            .in0(N__32713),
            .in1(N__29072),
            .in2(N__32860),
            .in3(N__33080),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_10_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_10_11_5 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_10_11_5  (
            .in0(N__33077),
            .in1(N__32815),
            .in2(N__29309),
            .in3(N__32712),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_11_6 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_10_11_6  (
            .in0(N__32715),
            .in1(N__28316),
            .in2(N__32862),
            .in3(N__33082),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_11_7 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_10_11_7  (
            .in0(N__33075),
            .in1(N__32810),
            .in2(N__28157),
            .in3(N__32709),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47937),
            .ce(N__32552),
            .sr(N__47323));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_10_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_10_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27575),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_12_4 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_12_4  (
            .in0(N__25460),
            .in1(_gnd_net_),
            .in2(N__25612),
            .in3(N__26397),
            .lcout(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_12_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_12_5  (
            .in0(N__26398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25605),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_10_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_10_12_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_10_12_6 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_10_12_6  (
            .in0(N__41279),
            .in1(N__35303),
            .in2(N__40730),
            .in3(N__40831),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47928),
            .ce(),
            .sr(N__47335));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_10_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_10_13_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_10_13_0  (
            .in0(N__25643),
            .in1(N__25503),
            .in2(N__26372),
            .in3(N__26337),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_10_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_10_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__30890),
            .in2(_gnd_net_),
            .in3(N__30801),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__25742),
            .in2(_gnd_net_),
            .in3(N__26771),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__30764),
            .in2(_gnd_net_),
            .in3(N__30843),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_10_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_10_13_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_10_13_4  (
            .in0(N__25770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26730),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__25642),
            .in2(_gnd_net_),
            .in3(N__26367),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_13_6  (
            .in0(N__26647),
            .in1(N__25836),
            .in2(N__25688),
            .in3(N__26599),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7  (
            .in0(N__26399),
            .in1(N__25641),
            .in2(N__25613),
            .in3(N__26368),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0  (
            .in0(N__26566),
            .in1(N__26194),
            .in2(N__26150),
            .in3(N__26538),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__25933),
            .in2(_gnd_net_),
            .in3(N__26689),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__26195),
            .in2(_gnd_net_),
            .in3(N__26539),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3  (
            .in0(N__25841),
            .in1(N__26146),
            .in2(N__26606),
            .in3(N__26565),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_14_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_14_4  (
            .in0(N__26304),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25890),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_14_5  (
            .in0(N__25505),
            .in1(N__25891),
            .in2(N__26342),
            .in3(N__26305),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__25504),
            .in2(_gnd_net_),
            .in3(N__26338),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_10_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_10_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_10_14_7  (
            .in0(N__25934),
            .in1(N__30805),
            .in2(N__26693),
            .in3(N__30886),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_10_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_10_15_0 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_10_15_0  (
            .in0(N__26878),
            .in1(_gnd_net_),
            .in2(N__26239),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_10_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_10_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_10_15_1  (
            .in0(N__26734),
            .in1(N__25932),
            .in2(N__25781),
            .in3(N__26688),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_15_2  (
            .in0(N__25892),
            .in1(N__26769),
            .in2(N__26309),
            .in3(N__25740),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_15_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__25837),
            .in2(_gnd_net_),
            .in3(N__26598),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_15_4 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_15_4  (
            .in0(N__25777),
            .in1(N__25741),
            .in2(N__26735),
            .in3(N__26770),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_15_5  (
            .in0(N__25989),
            .in1(N__26877),
            .in2(N__26921),
            .in3(N__26232),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_10_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_10_15_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_10_15_6  (
            .in0(N__26813),
            .in1(N__26069),
            .in2(N__30515),
            .in3(N__30465),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_15_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_15_7  (
            .in0(N__26068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26812),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_16_0 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_16_0  (
            .in0(N__26913),
            .in1(_gnd_net_),
            .in2(N__25994),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_16_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26024),
            .in3(N__26952),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_16_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26102),
            .in3(N__26841),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_10_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_10_16_3 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_10_16_3  (
            .in0(N__26842),
            .in1(N__26097),
            .in2(N__26885),
            .in3(N__26240),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_16_4 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_16_4  (
            .in0(N__26540),
            .in1(N__26019),
            .in2(N__26959),
            .in3(N__26188),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_16_5  (
            .in0(N__26140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26567),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_6  (
            .in0(N__26101),
            .in1(N__26067),
            .in2(N__26846),
            .in3(N__26806),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_7  (
            .in0(N__26023),
            .in1(N__25990),
            .in2(N__26960),
            .in3(N__26914),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_10_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_10_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__29735),
            .in2(N__29767),
            .in3(N__29763),
            .lcout(\current_shift_inst.un38_control_input_0 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_10_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_10_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__29723),
            .in2(_gnd_net_),
            .in3(N__26459),
            .lcout(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_10_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_10_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__29711),
            .in2(_gnd_net_),
            .in3(N__26423),
            .lcout(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_10_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_10_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__29834),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_10_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_10_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__29828),
            .in2(_gnd_net_),
            .in3(N__26375),
            .lcout(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_10_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_10_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__29822),
            .in2(_gnd_net_),
            .in3(N__26345),
            .lcout(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_10_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_10_17_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29816),
            .in3(N__26312),
            .lcout(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_10_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_10_17_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29807),
            .in3(N__26279),
            .lcout(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_10_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_10_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__29786),
            .in2(_gnd_net_),
            .in3(N__26738),
            .lcout(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_10_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_10_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__29780),
            .in2(_gnd_net_),
            .in3(N__26696),
            .lcout(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_10_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_10_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__29774),
            .in2(_gnd_net_),
            .in3(N__26657),
            .lcout(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_10_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_10_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__29888),
            .in2(_gnd_net_),
            .in3(N__26654),
            .lcout(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_10_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_10_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__29798),
            .in2(_gnd_net_),
            .in3(N__26651),
            .lcout(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_10_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_10_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__29717),
            .in2(_gnd_net_),
            .in3(N__26609),
            .lcout(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_10_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_10_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__29792),
            .in2(_gnd_net_),
            .in3(N__26570),
            .lcout(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_10_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_10_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__29882),
            .in2(_gnd_net_),
            .in3(N__26543),
            .lcout(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_10_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_10_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__29993),
            .in2(_gnd_net_),
            .in3(N__26513),
            .lcout(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_10_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_10_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__29870),
            .in2(_gnd_net_),
            .in3(N__26924),
            .lcout(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_10_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_10_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__29858),
            .in2(_gnd_net_),
            .in3(N__26888),
            .lcout(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_10_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_10_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__29876),
            .in2(_gnd_net_),
            .in3(N__26849),
            .lcout(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_10_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_10_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__29987),
            .in2(_gnd_net_),
            .in3(N__26816),
            .lcout(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_10_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_10_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__29846),
            .in2(_gnd_net_),
            .in3(N__26786),
            .lcout(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_10_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_10_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__29864),
            .in2(_gnd_net_),
            .in3(N__26783),
            .lcout(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_10_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_10_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__29840),
            .in2(_gnd_net_),
            .in3(N__26780),
            .lcout(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_10_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_10_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__29852),
            .in2(_gnd_net_),
            .in3(N__26777),
            .lcout(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_10_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_10_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__29978),
            .in2(_gnd_net_),
            .in3(N__26774),
            .lcout(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_10_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_10_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__29915),
            .in2(_gnd_net_),
            .in3(N__27179),
            .lcout(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_10_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_10_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__29897),
            .in2(_gnd_net_),
            .in3(N__27176),
            .lcout(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_10_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_10_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__29906),
            .in2(_gnd_net_),
            .in3(N__27173),
            .lcout(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_10_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_10_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__29924),
            .in2(_gnd_net_),
            .in3(N__27149),
            .lcout(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_29 ),
            .carryout(\current_shift_inst.un4_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_10_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__27134),
            .in2(_gnd_net_),
            .in3(N__27068),
            .lcout(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_10_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_10_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_10_20_7  (
            .in0(N__30697),
            .in1(N__27044),
            .in2(N__30655),
            .in3(N__27000),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_10_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_10_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_10_21_0  (
            .in0(N__27335),
            .in1(N__31086),
            .in2(_gnd_net_),
            .in3(N__26966),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_1_LC_10_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_10_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_10_21_1  (
            .in0(N__27330),
            .in1(N__31047),
            .in2(_gnd_net_),
            .in3(N__26963),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_2_LC_10_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_10_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_10_21_2  (
            .in0(N__27336),
            .in1(N__31017),
            .in2(_gnd_net_),
            .in3(N__27206),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_3_LC_10_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_10_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_10_21_3  (
            .in0(N__27331),
            .in1(N__30987),
            .in2(_gnd_net_),
            .in3(N__27203),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_4_LC_10_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_10_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_10_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_10_21_4  (
            .in0(N__27337),
            .in1(N__30946),
            .in2(_gnd_net_),
            .in3(N__27200),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_5_LC_10_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_10_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_10_21_5  (
            .in0(N__27332),
            .in1(N__30910),
            .in2(_gnd_net_),
            .in3(N__27197),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_6_LC_10_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_10_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_10_21_6  (
            .in0(N__27334),
            .in1(N__31615),
            .in2(_gnd_net_),
            .in3(N__27194),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_7_LC_10_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_10_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_10_21_7  (
            .in0(N__27333),
            .in1(N__31585),
            .in2(_gnd_net_),
            .in3(N__27191),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__47877),
            .ce(N__27517),
            .sr(N__47399));
    defparam \current_shift_inst.timer_s1.counter_8_LC_10_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_10_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_10_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_10_22_0  (
            .in0(N__27341),
            .in1(N__31551),
            .in2(_gnd_net_),
            .in3(N__27188),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_9_LC_10_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_10_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_10_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_10_22_1  (
            .in0(N__27345),
            .in1(N__31509),
            .in2(_gnd_net_),
            .in3(N__27185),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_10_LC_10_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_10_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_10_22_2  (
            .in0(N__27338),
            .in1(N__31470),
            .in2(_gnd_net_),
            .in3(N__27182),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_11_LC_10_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_10_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_10_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_10_22_3  (
            .in0(N__27342),
            .in1(N__31434),
            .in2(_gnd_net_),
            .in3(N__27236),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_12_LC_10_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_10_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_10_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_10_22_4  (
            .in0(N__27339),
            .in1(N__31396),
            .in2(_gnd_net_),
            .in3(N__27233),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_13_LC_10_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_10_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_10_22_5  (
            .in0(N__27343),
            .in1(N__31900),
            .in2(_gnd_net_),
            .in3(N__27230),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_14_LC_10_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_10_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_10_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_10_22_6  (
            .in0(N__27340),
            .in1(N__31864),
            .in2(_gnd_net_),
            .in3(N__27227),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_15_LC_10_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_10_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_10_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_10_22_7  (
            .in0(N__27344),
            .in1(N__31828),
            .in2(_gnd_net_),
            .in3(N__27224),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__47870),
            .ce(N__27518),
            .sr(N__47403));
    defparam \current_shift_inst.timer_s1.counter_16_LC_10_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_10_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_10_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_10_23_0  (
            .in0(N__27350),
            .in1(N__31797),
            .in2(_gnd_net_),
            .in3(N__27221),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_17_LC_10_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_10_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_10_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_10_23_1  (
            .in0(N__27346),
            .in1(N__31758),
            .in2(_gnd_net_),
            .in3(N__27218),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_18_LC_10_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_10_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_10_23_2  (
            .in0(N__27351),
            .in1(N__31719),
            .in2(_gnd_net_),
            .in3(N__27215),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_19_LC_10_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_10_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_10_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_10_23_3  (
            .in0(N__27347),
            .in1(N__31683),
            .in2(_gnd_net_),
            .in3(N__27212),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_20_LC_10_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_10_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_10_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_10_23_4  (
            .in0(N__27352),
            .in1(N__31648),
            .in2(_gnd_net_),
            .in3(N__27209),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_21_LC_10_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_10_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_10_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_10_23_5  (
            .in0(N__27348),
            .in1(N__32239),
            .in2(_gnd_net_),
            .in3(N__27383),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_22_LC_10_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_10_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_10_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_10_23_6  (
            .in0(N__27353),
            .in1(N__32203),
            .in2(_gnd_net_),
            .in3(N__27380),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_23_LC_10_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_10_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_10_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_10_23_7  (
            .in0(N__27349),
            .in1(N__32167),
            .in2(_gnd_net_),
            .in3(N__27377),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__47864),
            .ce(N__27507),
            .sr(N__47406));
    defparam \current_shift_inst.timer_s1.counter_24_LC_10_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_10_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_10_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_10_24_0  (
            .in0(N__27354),
            .in1(N__32136),
            .in2(_gnd_net_),
            .in3(N__27374),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__47859),
            .ce(N__27506),
            .sr(N__47410));
    defparam \current_shift_inst.timer_s1.counter_25_LC_10_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_10_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_10_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_10_24_1  (
            .in0(N__27358),
            .in1(N__32097),
            .in2(_gnd_net_),
            .in3(N__27371),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__47859),
            .ce(N__27506),
            .sr(N__47410));
    defparam \current_shift_inst.timer_s1.counter_26_LC_10_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_10_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_10_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_10_24_2  (
            .in0(N__27355),
            .in1(N__32040),
            .in2(_gnd_net_),
            .in3(N__27368),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__47859),
            .ce(N__27506),
            .sr(N__47410));
    defparam \current_shift_inst.timer_s1.counter_27_LC_10_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_10_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_10_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_10_24_3  (
            .in0(N__27359),
            .in1(N__31986),
            .in2(_gnd_net_),
            .in3(N__27365),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__47859),
            .ce(N__27506),
            .sr(N__47410));
    defparam \current_shift_inst.timer_s1.counter_28_LC_10_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_10_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_10_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_10_24_4  (
            .in0(N__27356),
            .in1(N__32062),
            .in2(_gnd_net_),
            .in3(N__27362),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__47859),
            .ce(N__27506),
            .sr(N__47410));
    defparam \current_shift_inst.timer_s1.counter_29_LC_10_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_10_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_10_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_10_24_5  (
            .in0(N__32008),
            .in1(N__27357),
            .in2(_gnd_net_),
            .in3(N__27239),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47859),
            .ce(N__27506),
            .sr(N__47410));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_10_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_10_25_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_10_25_4  (
            .in0(N__27601),
            .in1(N__27567),
            .in2(_gnd_net_),
            .in3(N__27540),
            .lcout(\current_shift_inst.timer_s1.N_192_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_phase_LC_10_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_phase_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_phase_LC_10_25_6 .LUT_INIT=16'b1011101110100000;
    LogicCell40 \current_shift_inst.stop_timer_phase_LC_10_25_6  (
            .in0(N__30285),
            .in1(N__30233),
            .in2(N__32305),
            .in3(N__27451),
            .lcout(\current_shift_inst.stop_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47853),
            .ce(N__35836),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_10_26_3.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_10_26_3.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_10_26_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_10_26_3 (
            .in0(N__47460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_10_26_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_10_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIC90O_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(N__27470),
            .in2(_gnd_net_),
            .in3(N__27446),
            .lcout(\current_shift_inst.timer_phase.N_188_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_11_5_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_11_5_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_11_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27410),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47973),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_11_6_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_11_6_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_11_6_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_11_6_2 (
            .in0(N__27398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47964),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_11_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_11_9_0 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_11_9_0  (
            .in0(N__32896),
            .in1(N__33007),
            .in2(N__28766),
            .in3(N__32691),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47947),
            .ce(N__32551),
            .sr(N__47304));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_9_1 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_11_9_1  (
            .in0(N__32694),
            .in1(N__33010),
            .in2(N__27626),
            .in3(N__32899),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47947),
            .ce(N__32551),
            .sr(N__47304));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_11_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_11_9_3 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_11_9_3  (
            .in0(N__32693),
            .in1(N__33009),
            .in2(N__27704),
            .in3(N__32898),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47947),
            .ce(N__32551),
            .sr(N__47304));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_9_4 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_11_9_4  (
            .in0(N__32897),
            .in1(N__33008),
            .in2(N__29654),
            .in3(N__32692),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47947),
            .ce(N__32551),
            .sr(N__47304));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_11_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_11_9_5 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_11_9_5  (
            .in0(N__30125),
            .in1(N__32895),
            .in2(N__27938),
            .in3(N__30082),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47947),
            .ce(N__32551),
            .sr(N__47304));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__27984),
            .in2(N__27964),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un1_integrator_axb_0 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__27918),
            .in2(N__27899),
            .in3(N__27866),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__30024),
            .in2(N__27863),
            .in3(N__27839),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__27832),
            .in2(N__27803),
            .in3(N__27764),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__27744),
            .in2(N__27728),
            .in3(N__27695),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__27677),
            .in2(N__27655),
            .in3(N__27617),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__28505),
            .in2(N__28484),
            .in3(N__28451),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__28423),
            .in2(N__28411),
            .in3(N__28376),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__28361),
            .in2(N__28340),
            .in3(N__28307),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__28286),
            .in2(N__28261),
            .in3(N__28223),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__28195),
            .in2(N__28183),
            .in3(N__28148),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__28134),
            .in2(N__28109),
            .in3(N__28073),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__28050),
            .in2(N__28034),
            .in3(N__27995),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__29045),
            .in2(N__29024),
            .in3(N__28988),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__28980),
            .in2(N__28955),
            .in3(N__28913),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__28902),
            .in2(N__28877),
            .in3(N__28844),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__28826),
            .in2(N__28793),
            .in3(N__28754),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__28743),
            .in2(N__28712),
            .in3(N__28673),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__28663),
            .in2(N__28634),
            .in3(N__28595),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__28590),
            .in2(N__28556),
            .in3(N__28520),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__29446),
            .in2(N__29422),
            .in3(N__29369),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__29356),
            .in2(N__29336),
            .in3(N__29300),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__29291),
            .in2(N__29258),
            .in3(N__29225),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__29218),
            .in2(N__29186),
            .in3(N__29150),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__30403),
            .in2(N__29147),
            .in3(N__29120),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__30349),
            .in2(N__29506),
            .in3(N__29117),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__29491),
            .in2(N__29107),
            .in3(N__29063),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__32597),
            .in2(N__29507),
            .in3(N__29060),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__29495),
            .in2(N__29704),
            .in3(N__29639),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__29632),
            .in2(N__29508),
            .in3(N__29579),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__29499),
            .in2(N__29575),
            .in3(N__29513),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_13_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_13_7  (
            .in0(N__33041),
            .in1(_gnd_net_),
            .in2(N__29509),
            .in3(N__29453),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_14_0 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_11_14_0  (
            .in0(N__34844),
            .in1(N__34768),
            .in2(N__39728),
            .in3(N__34856),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47910),
            .ce(N__33561),
            .sr(N__47344));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_14_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_11_14_7  (
            .in0(N__34963),
            .in1(N__40529),
            .in2(_gnd_net_),
            .in3(N__35143),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47910),
            .ce(N__33561),
            .sr(N__47344));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_c_0_LC_11_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_c_0_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_c_0_LC_11_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_c_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__40510),
            .in2(_gnd_net_),
            .in3(N__33142),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_15_2 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_11_15_2  (
            .in0(N__40511),
            .in1(N__35604),
            .in2(N__29450),
            .in3(N__34816),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47904),
            .ce(N__33565),
            .sr(N__47354));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31099),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47897),
            .ce(N__31958),
            .sr(N__47362));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31060),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47897),
            .ce(N__31958),
            .sr(N__47362));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31927),
            .lcout(\current_shift_inst.elapsed_time_ns_1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47897),
            .ce(N__31958),
            .sr(N__47362));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_17_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_11_17_2  (
            .in0(N__34988),
            .in1(_gnd_net_),
            .in2(N__40558),
            .in3(N__34517),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47891),
            .ce(N__33556),
            .sr(N__47372));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_17_3 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_17_3  (
            .in0(N__35057),
            .in1(N__40547),
            .in2(_gnd_net_),
            .in3(N__34987),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47891),
            .ce(N__33556),
            .sr(N__47372));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_4  (
            .in0(N__40546),
            .in1(N__36800),
            .in2(_gnd_net_),
            .in3(N__35228),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47891),
            .ce(N__33556),
            .sr(N__47372));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29741),
            .lcout(\current_shift_inst.un4_control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29729),
            .lcout(\current_shift_inst.un4_control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_11_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_11_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31415),
            .lcout(\current_shift_inst.un4_control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31067),
            .lcout(\current_shift_inst.un4_control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31028),
            .lcout(\current_shift_inst.un4_control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30998),
            .lcout(\current_shift_inst.un4_control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30968),
            .lcout(\current_shift_inst.un4_control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30932),
            .lcout(\current_shift_inst.un4_control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30896),
            .lcout(\current_shift_inst.un4_control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_11_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_11_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31451),
            .lcout(\current_shift_inst.un4_control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31382),
            .lcout(\current_shift_inst.un4_control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31601),
            .lcout(\current_shift_inst.un4_control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_11_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_11_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31571),
            .lcout(\current_shift_inst.un4_control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_11_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_11_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31529),
            .lcout(\current_shift_inst.un4_control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31487),
            .lcout(\current_shift_inst.un4_control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_11_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_11_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31886),
            .lcout(\current_shift_inst.un4_control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_11_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_11_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31736),
            .lcout(\current_shift_inst.un4_control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_11_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_11_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31814),
            .lcout(\current_shift_inst.un4_control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31634),
            .lcout(\current_shift_inst.un4_control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_11_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_11_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31775),
            .lcout(\current_shift_inst.un4_control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32189),
            .lcout(\current_shift_inst.un4_control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_11_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_11_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31664),
            .lcout(\current_shift_inst.un4_control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_11_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_11_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32225),
            .lcout(\current_shift_inst.un4_control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31850),
            .lcout(\current_shift_inst.un4_control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_11_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_11_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31700),
            .lcout(\current_shift_inst.un4_control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32153),
            .lcout(\current_shift_inst.un4_control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_11_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_11_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_i_31_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29968),
            .lcout(\current_shift_inst.z_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31967),
            .lcout(\current_shift_inst.un4_control_input_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_11_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_11_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32114),
            .lcout(\current_shift_inst.un4_control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_11_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_11_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32021),
            .lcout(\current_shift_inst.un4_control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32075),
            .lcout(\current_shift_inst.un4_control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_rise_LC_11_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.S1_rise_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_rise_LC_11_24_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S1_rise_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__30314),
            .in2(_gnd_net_),
            .in3(N__30301),
            .lcout(\current_shift_inst.S1_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47854),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync0_LC_11_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync0_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync0_LC_11_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync0_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32317),
            .lcout(\current_shift_inst.S1_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47854),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync_prev_LC_11_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync_prev_LC_11_24_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync_prev_LC_11_24_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S1_sync_prev_LC_11_24_4  (
            .in0(N__30302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S1_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47854),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync1_LC_11_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync1_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync1_LC_11_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync1_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30308),
            .lcout(\current_shift_inst.S1_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47854),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.phase_valid_LC_11_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_LC_11_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.phase_valid_LC_11_25_7 .LUT_INIT=16'b1100100011101010;
    LogicCell40 \current_shift_inst.phase_valid_LC_11_25_7  (
            .in0(N__30184),
            .in1(N__30293),
            .in2(N__32292),
            .in3(N__30232),
            .lcout(\current_shift_inst.phase_validZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__47411));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_12_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30137),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47962),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_5_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_5_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_5_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_12_5_7 (
            .in0(N__30152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47962),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_12_7_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_12_7_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_12_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_12_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30131),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47954),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_12_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_12_9_4 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_12_9_4  (
            .in0(N__30124),
            .in1(N__32909),
            .in2(N__30086),
            .in3(N__30047),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47936),
            .ce(N__32554),
            .sr(N__47297));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_12_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_12_10_7 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_12_10_7  (
            .in0(N__33003),
            .in1(N__32900),
            .in2(N__30008),
            .in3(N__32720),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47927),
            .ce(N__32555),
            .sr(N__47305));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_1 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_1  (
            .in0(N__33004),
            .in1(N__32891),
            .in2(N__30419),
            .in3(N__32721),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47921),
            .ce(N__32530),
            .sr(N__47312));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_12_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_12_11_2 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_12_11_2  (
            .in0(N__32722),
            .in1(N__30365),
            .in2(N__32907),
            .in3(N__33005),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47921),
            .ce(N__32530),
            .sr(N__47312));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_12_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_12_0  (
            .in0(N__39958),
            .in1(N__40232),
            .in2(N__40127),
            .in3(N__37220),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47914),
            .ce(),
            .sr(N__47318));
    defparam \phase_controller_inst1.stoper_hc.un1_m5_i_1_LC_12_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m5_i_1_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m5_i_1_LC_12_12_4 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m5_i_1_LC_12_12_4  (
            .in0(N__35039),
            .in1(N__33119),
            .in2(N__36419),
            .in3(N__33113),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_m5_iZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m5_i_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m5_i_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m5_i_LC_12_12_5 .LUT_INIT=16'b1111101110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m5_i_LC_12_12_5  (
            .in0(N__35180),
            .in1(N__32333),
            .in2(N__30320),
            .in3(N__39724),
            .lcout(\phase_controller_inst1.stoper_hc.un1_N_4 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_12_6 .LUT_INIT=16'b0011111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__34893),
            .in2(N__30317),
            .in3(N__33130),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_12_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_12_13_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_12_13_0  (
            .in0(N__40519),
            .in1(N__34648),
            .in2(_gnd_net_),
            .in3(N__34948),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47909),
            .ce(N__33540),
            .sr(N__47324));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1  (
            .in0(N__35448),
            .in1(N__35542),
            .in2(N__34607),
            .in3(N__40524),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47909),
            .ce(N__33540),
            .sr(N__47324));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_13_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_12_13_2  (
            .in0(N__35541),
            .in1(N__34561),
            .in2(N__40552),
            .in3(N__35450),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47909),
            .ce(N__33540),
            .sr(N__47324));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_13_3 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_12_13_3  (
            .in0(N__35449),
            .in1(N__35543),
            .in2(N__35278),
            .in3(N__40525),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47909),
            .ce(N__33540),
            .sr(N__47324));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_13_4 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_12_13_4  (
            .in0(N__35540),
            .in1(N__35311),
            .in2(N__40551),
            .in3(N__35447),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47909),
            .ce(N__33540),
            .sr(N__47324));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_12_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_12_13_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_12_13_5  (
            .in0(N__34949),
            .in1(N__40520),
            .in2(_gnd_net_),
            .in3(N__39766),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47909),
            .ce(N__33540),
            .sr(N__47324));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_14_0 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_14_0  (
            .in0(N__40062),
            .in1(N__40200),
            .in2(N__36926),
            .in3(N__39936),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47903),
            .ce(),
            .sr(N__47336));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_1  (
            .in0(N__40199),
            .in1(N__40065),
            .in2(N__39961),
            .in3(N__37166),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47903),
            .ce(),
            .sr(N__47336));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2  (
            .in0(N__40061),
            .in1(N__39937),
            .in2(N__37136),
            .in3(N__40201),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47903),
            .ce(),
            .sr(N__47336));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_14_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_14_3  (
            .in0(N__40197),
            .in1(N__40063),
            .in2(N__39959),
            .in3(N__33440),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47903),
            .ce(),
            .sr(N__47336));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_14_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_14_7  (
            .in0(N__40198),
            .in1(N__40064),
            .in2(N__39960),
            .in3(N__36890),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47903),
            .ce(),
            .sr(N__47336));
    defparam \phase_controller_inst1.state_3_LC_12_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_15_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_15_0  (
            .in0(N__33851),
            .in1(N__34410),
            .in2(N__34450),
            .in3(N__33749),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47896),
            .ce(),
            .sr(N__47345));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_12_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_12_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__34321),
            .in2(_gnd_net_),
            .in3(N__34285),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_12_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_12_16_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__37774),
            .in2(_gnd_net_),
            .in3(N__38047),
            .lcout(\phase_controller_slave.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_12_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_12_16_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_12_16_1  (
            .in0(N__38048),
            .in1(N__37973),
            .in2(_gnd_net_),
            .in3(N__37780),
            .lcout(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_12_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_12_16_6 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_12_16_6  (
            .in0(N__34904),
            .in1(N__33146),
            .in2(N__40509),
            .in3(N__34873),
            .lcout(\phase_controller_inst1.stoper_hc.un1_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_12_17_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_12_17_0  (
            .in0(N__30885),
            .in1(N__30844),
            .in2(N__30809),
            .in3(N__30763),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_12_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_12_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__33950),
            .in2(_gnd_net_),
            .in3(N__33987),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_17_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__31283),
            .in2(_gnd_net_),
            .in3(N__31188),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_12_17_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_12_17_4  (
            .in0(N__31373),
            .in1(N__30698),
            .in2(N__31337),
            .in3(N__30654),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_12_17_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_12_17_5  (
            .in0(N__30508),
            .in1(N__30602),
            .in2(N__30470),
            .in3(N__30561),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_12_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_12_17_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__30507),
            .in2(_gnd_net_),
            .in3(N__30466),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_12_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__31372),
            .in2(_gnd_net_),
            .in3(N__31332),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_12_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_12_18_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_12_18_5  (
            .in0(N__31282),
            .in1(N__31230),
            .in2(N__31193),
            .in3(N__31145),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__31018),
            .in2(N__31100),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__30988),
            .in2(N__31061),
            .in3(N__31022),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__31019),
            .in2(N__30958),
            .in3(N__30992),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__30989),
            .in2(N__30922),
            .in3(N__30962),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__31621),
            .in2(N__30959),
            .in3(N__30926),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__31591),
            .in2(N__30923),
            .in3(N__31625),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__31622),
            .in2(N__31562),
            .in3(N__31595),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__31592),
            .in2(N__31520),
            .in3(N__31565),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47876),
            .ce(N__31957),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__31561),
            .in2(N__31477),
            .in3(N__31523),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__31519),
            .in2(N__31441),
            .in3(N__31481),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__31402),
            .in2(N__31478),
            .in3(N__31445),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__31906),
            .in2(N__31442),
            .in3(N__31406),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__31403),
            .in2(N__31876),
            .in3(N__31376),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__31907),
            .in2(N__31840),
            .in3(N__31880),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__31804),
            .in2(N__31877),
            .in3(N__31844),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__31765),
            .in2(N__31841),
            .in3(N__31808),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47869),
            .ce(N__31956),
            .sr(N__47383));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__31805),
            .in2(N__31726),
            .in3(N__31769),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__31766),
            .in2(N__31690),
            .in3(N__31730),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__31654),
            .in2(N__31727),
            .in3(N__31694),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__32245),
            .in2(N__31691),
            .in3(N__31658),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__31655),
            .in2(N__32215),
            .in3(N__31628),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__32246),
            .in2(N__32179),
            .in3(N__32219),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__32143),
            .in2(N__32216),
            .in3(N__32183),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__32104),
            .in2(N__32180),
            .in3(N__32147),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47863),
            .ce(N__31955),
            .sr(N__47391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__32144),
            .in2(N__32047),
            .in3(N__32108),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47858),
            .ce(N__31954),
            .sr(N__47395));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__32105),
            .in2(N__31993),
            .in3(N__32069),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47858),
            .ce(N__31954),
            .sr(N__47395));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__32066),
            .in2(N__32048),
            .in3(N__32015),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47858),
            .ce(N__31954),
            .sr(N__47395));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__32012),
            .in2(N__31994),
            .in3(N__31961),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47858),
            .ce(N__31954),
            .sr(N__47395));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31934),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_23_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_23_2  (
            .in0(N__36102),
            .in1(N__36054),
            .in2(_gnd_net_),
            .in3(N__36279),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_12_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_12_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_12_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34457),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_25_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_12_25_0  (
            .in0(N__48338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47849),
            .ce(N__43111),
            .sr(N__47407));
    defparam \current_shift_inst.S3_rise_LC_12_26_0 .C_ON=1'b0;
    defparam \current_shift_inst.S3_rise_LC_12_26_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_rise_LC_12_26_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S3_rise_LC_12_26_0  (
            .in0(_gnd_net_),
            .in1(N__32267),
            .in2(_gnd_net_),
            .in3(N__32254),
            .lcout(\current_shift_inst.S3_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47848),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync0_LC_12_26_1 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync0_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync0_LC_12_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync0_LC_12_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33895),
            .lcout(\current_shift_inst.S3_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47848),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync_prev_LC_12_26_2 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync_prev_LC_12_26_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync_prev_LC_12_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync_prev_LC_12_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32255),
            .lcout(\current_shift_inst.S3_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47848),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_12_26_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_12_26_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_12_26_4  (
            .in0(_gnd_net_),
            .in1(N__36017),
            .in2(_gnd_net_),
            .in3(N__36278),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync1_LC_12_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync1_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync1_LC_12_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync1_LC_12_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32261),
            .lcout(\current_shift_inst.S3_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47848),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_13_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_13_6_0 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_13_6_0  (
            .in0(N__36574),
            .in1(N__36552),
            .in2(_gnd_net_),
            .in3(N__36452),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47965),
            .ce(N__35897),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_13_7_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_13_7_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_13_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_13_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33095),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47957),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_8_7  (
            .in0(N__34641),
            .in1(N__36403),
            .in2(N__35350),
            .in3(N__35046),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_9_1 .LUT_INIT=16'b1111101101110011;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_13_9_1  (
            .in0(N__40718),
            .in1(N__36698),
            .in2(N__34807),
            .in3(N__44228),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47948),
            .ce(),
            .sr(N__47292));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_13_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_13_9_5 .LUT_INIT=16'b1111101101110011;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_13_9_5  (
            .in0(N__40719),
            .in1(N__36699),
            .in2(N__34732),
            .in3(N__44285),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47948),
            .ce(),
            .sr(N__47292));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_9_6 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_13_9_6  (
            .in0(N__35131),
            .in1(N__40720),
            .in2(N__41396),
            .in3(N__40853),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47948),
            .ce(),
            .sr(N__47292));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_9_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_13_9_7  (
            .in0(N__40717),
            .in1(N__35176),
            .in2(N__42016),
            .in3(N__36700),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47948),
            .ce(),
            .sr(N__47292));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_13_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_13_10_4 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_13_10_4  (
            .in0(N__33006),
            .in1(N__32908),
            .in2(N__32738),
            .in3(N__32723),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47938),
            .ce(N__32561),
            .sr(N__47298));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_13_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_13_11_0  (
            .in0(N__34673),
            .in1(N__34636),
            .in2(N__35368),
            .in3(N__35136),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_13_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_13_11_2 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_13_11_2  (
            .in0(N__34640),
            .in1(N__40722),
            .in2(N__41495),
            .in3(N__40844),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47929),
            .ce(),
            .sr(N__47306));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_13_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_13_11_4 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_13_11_4  (
            .in0(N__35045),
            .in1(N__40723),
            .in2(N__44021),
            .in3(N__40845),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47929),
            .ce(),
            .sr(N__47306));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_13_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_13_11_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_13_11_6  (
            .in0(N__33155),
            .in1(N__34208),
            .in2(N__39723),
            .in3(N__34220),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_13_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_13_12_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_13_12_0  (
            .in0(N__36823),
            .in1(N__36724),
            .in2(N__36767),
            .in3(N__35213),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_13_12_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_13_12_1  (
            .in0(N__35489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34556),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_LC_13_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_LC_13_12_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_LC_13_12_2  (
            .in0(N__39591),
            .in1(N__34201),
            .in2(N__35274),
            .in3(N__34219),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_13_12_3 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_13_12_3  (
            .in0(N__34202),
            .in1(N__34193),
            .in2(_gnd_net_),
            .in3(N__35267),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_13_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_13_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_LC_13_12_4  (
            .in0(N__36792),
            .in1(N__33107),
            .in2(N__33101),
            .in3(N__35214),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlt31 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlt31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_12_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33098),
            .in3(N__40461),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_12_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_12_6  (
            .in0(N__39938),
            .in1(N__40006),
            .in2(_gnd_net_),
            .in3(N__40202),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_13_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__42785),
            .in2(_gnd_net_),
            .in3(N__42989),
            .lcout(\phase_controller_slave.start_timer_hc_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__33293),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__33266),
            .in2(N__33275),
            .in3(N__37026),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__33251),
            .in2(N__33260),
            .in3(N__37009),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__33236),
            .in2(N__33245),
            .in3(N__36964),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__33230),
            .in2(N__33224),
            .in3(N__36937),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__33200),
            .in2(N__33215),
            .in3(N__36901),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__33179),
            .in2(N__33194),
            .in3(N__36874),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__33161),
            .in2(N__33173),
            .in3(N__37231),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__33422),
            .in2(N__33434),
            .in3(N__37204),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__33392),
            .in2(N__33416),
            .in3(N__37177),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__33368),
            .in2(N__33386),
            .in3(N__40301),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__33350),
            .in2(N__33362),
            .in3(N__37147),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__33344),
            .in2(N__33599),
            .in3(N__37120),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_14_5  (
            .in0(N__40280),
            .in1(N__33323),
            .in2(N__33338),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__33305),
            .in2(N__33317),
            .in3(N__37096),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__33299),
            .in2(N__33614),
            .in3(N__40259),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__33482),
            .in2(N__33494),
            .in3(N__37373),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__33476),
            .in2(N__33587),
            .in3(N__37346),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_15_2  (
            .in0(N__37321),
            .in1(N__33470),
            .in2(N__33578),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__33449),
            .in2(N__33464),
            .in3(N__39836),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33443),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_15_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_15_5  (
            .in0(N__40060),
            .in1(N__39923),
            .in2(_gnd_net_),
            .in3(N__40193),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_13_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_13_15_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_13_15_7  (
            .in0(N__34322),
            .in1(N__37030),
            .in2(_gnd_net_),
            .in3(N__34286),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_16_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_13_16_0  (
            .in0(N__35414),
            .in1(N__35597),
            .in2(N__40536),
            .in3(N__35499),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47898),
            .ce(N__33557),
            .sr(N__47346));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_16_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_13_16_1  (
            .in0(N__35594),
            .in1(N__40488),
            .in2(N__35194),
            .in3(N__35412),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47898),
            .ce(N__33557),
            .sr(N__47346));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_16_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_13_16_3  (
            .in0(N__35369),
            .in1(N__40487),
            .in2(_gnd_net_),
            .in3(N__34992),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47898),
            .ce(N__33557),
            .sr(N__47346));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_13_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_13_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_13_16_4 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_13_16_4  (
            .in0(N__40489),
            .in1(N__35595),
            .in2(N__34742),
            .in3(N__34775),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47898),
            .ce(N__33557),
            .sr(N__47346));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_13_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_13_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_13_16_6 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_13_16_6  (
            .in0(N__35413),
            .in1(N__35596),
            .in2(N__40535),
            .in3(N__35096),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47898),
            .ce(N__33557),
            .sr(N__47346));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_17_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_17_0  (
            .in0(N__39915),
            .in1(N__40184),
            .in2(N__40100),
            .in3(N__34294),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_13_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_13_17_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_13_17_1  (
            .in0(N__34295),
            .in1(N__40066),
            .in2(N__40229),
            .in3(N__39916),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_17_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_17_2  (
            .in0(N__36065),
            .in1(N__36245),
            .in2(N__36204),
            .in3(N__39219),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_17_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_17_4  (
            .in0(N__43519),
            .in1(N__43032),
            .in2(N__43733),
            .in3(N__43790),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_17_5 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_17_5  (
            .in0(N__43033),
            .in1(N__43728),
            .in2(N__43833),
            .in3(N__43520),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_17_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_17_6  (
            .in0(N__37792),
            .in1(N__37974),
            .in2(N__38104),
            .in3(N__38698),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_17_7 .LUT_INIT=16'b0011000001000100;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_17_7  (
            .in0(N__38699),
            .in1(N__38062),
            .in2(N__38008),
            .in3(N__37793),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47892),
            .ce(N__35887),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_13_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_13_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_13_18_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_13_18_0  (
            .in0(N__37791),
            .in1(N__38058),
            .in2(N__37972),
            .in3(N__35630),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47885),
            .ce(),
            .sr(N__47363));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_13_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_13_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_13_18_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_13_18_3  (
            .in0(N__33778),
            .in1(N__38189),
            .in2(N__33794),
            .in3(N__38697),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47885),
            .ce(),
            .sr(N__47363));
    defparam \phase_controller_slave.state_0_LC_13_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_13_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_13_18_4 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_slave.state_0_LC_13_18_4  (
            .in0(N__33761),
            .in1(N__33994),
            .in2(N__33779),
            .in3(N__33945),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47885),
            .ce(),
            .sr(N__47363));
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_13_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_13_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_RNIVDE2_0_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__33774),
            .in2(_gnd_net_),
            .in3(N__33760),
            .lcout(\phase_controller_slave.state_RNIVDE2Z0Z_0 ),
            .ltout(\phase_controller_slave.state_RNIVDE2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_3_LC_13_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_13_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_13_18_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_slave.state_3_LC_13_18_6  (
            .in0(N__42813),
            .in1(N__42861),
            .in2(N__33752),
            .in3(N__33742),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47885),
            .ce(),
            .sr(N__47363));
    defparam \phase_controller_slave.state_ns_i_a2_1_LC_13_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.state_ns_i_a2_1_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_ns_i_a2_1_LC_13_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_ns_i_a2_1_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__33718),
            .in2(_gnd_net_),
            .in3(N__42891),
            .lcout(state_ns_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_13_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_19_2 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_19_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_19_2  (
            .in0(N__33729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42892),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47882),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_slave.S2_LC_13_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_13_19_3 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \phase_controller_slave.S2_LC_13_19_3  (
            .in0(N__33625),
            .in1(N__42812),
            .in2(N__33872),
            .in3(N__33941),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47882),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_slave.state_1_LC_13_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_13_19_4 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_slave.state_1_LC_13_19_4  (
            .in0(N__33995),
            .in1(N__42781),
            .in2(N__33949),
            .in3(N__42988),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47882),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_slave.start_timer_tr_LC_13_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_13_19_5 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_13_19_5  (
            .in0(N__42893),
            .in1(N__37921),
            .in2(N__33920),
            .in3(N__33908),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47882),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_slave.S1_LC_13_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_13_20_4 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \phase_controller_slave.S1_LC_13_20_4  (
            .in0(N__42817),
            .in1(_gnd_net_),
            .in2(N__33871),
            .in3(N__33883),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47878),
            .ce(),
            .sr(N__47378));
    defparam \phase_controller_inst1.T23_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_13_20_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \phase_controller_inst1.T23_LC_13_20_7  (
            .in0(N__34142),
            .in1(N__33864),
            .in2(_gnd_net_),
            .in3(N__34453),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47878),
            .ce(),
            .sr(N__47378));
    defparam \phase_controller_inst1.start_timer_tr_LC_13_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_22_0 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_13_22_0  (
            .in0(N__33844),
            .in1(N__33824),
            .in2(N__36176),
            .in3(N__42904),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47865),
            .ce(),
            .sr(N__47392));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_13_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_13_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__33813),
            .in2(_gnd_net_),
            .in3(N__33802),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_23_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_23_3  (
            .in0(N__33817),
            .in1(N__34252),
            .in2(N__33833),
            .in3(N__39220),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47860),
            .ce(),
            .sr(N__47396));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__34136),
            .in2(_gnd_net_),
            .in3(N__34177),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_13_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_13_23_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst1.state_0_LC_13_23_5  (
            .in0(N__33803),
            .in1(N__34178),
            .in2(N__33818),
            .in3(N__34140),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47860),
            .ce(),
            .sr(N__47396));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_23_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_23_6  (
            .in0(N__36060),
            .in1(N__36255),
            .in2(N__36180),
            .in3(N__34037),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47860),
            .ce(),
            .sr(N__47396));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_13_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_13_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__34091),
            .in2(N__38620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_13_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_13_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__38591),
            .in2(_gnd_net_),
            .in3(N__34019),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_13_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_13_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__34082),
            .in2(N__38570),
            .in3(N__34016),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_13_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_13_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__38909),
            .in2(_gnd_net_),
            .in3(N__34013),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_13_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_13_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__38891),
            .in2(_gnd_net_),
            .in3(N__34010),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_13_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_13_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__38873),
            .in2(_gnd_net_),
            .in3(N__34007),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_13_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_13_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__38852),
            .in2(_gnd_net_),
            .in3(N__34004),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_13_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_13_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__38834),
            .in2(_gnd_net_),
            .in3(N__34001),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_13_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_13_25_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38816),
            .in3(N__33998),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_13_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_13_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__38789),
            .in2(_gnd_net_),
            .in3(N__34055),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_13_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_13_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(N__39074),
            .in2(_gnd_net_),
            .in3(N__34052),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_13_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_13_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_13_25_3  (
            .in0(_gnd_net_),
            .in1(N__39056),
            .in2(_gnd_net_),
            .in3(N__34049),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_13_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_13_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(N__39038),
            .in2(_gnd_net_),
            .in3(N__34046),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_13_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_13_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(N__39020),
            .in2(_gnd_net_),
            .in3(N__34043),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_13_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_13_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(N__39002),
            .in2(_gnd_net_),
            .in3(N__34040),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_13_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_13_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_13_25_7  (
            .in0(_gnd_net_),
            .in1(N__38968),
            .in2(_gnd_net_),
            .in3(N__34028),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_13_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_13_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__38945),
            .in2(_gnd_net_),
            .in3(N__34025),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_13_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_13_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__38927),
            .in2(_gnd_net_),
            .in3(N__34022),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_13_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_13_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__39242),
            .in2(_gnd_net_),
            .in3(N__34094),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_26_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__34238),
            .in2(_gnd_net_),
            .in3(N__39205),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_13_26_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_13_26_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_13_26_7  (
            .in0(N__39206),
            .in1(_gnd_net_),
            .in2(N__34248),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_30_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_30_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34141),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(),
            .sr(N__47421));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_6  (
            .in0(N__39104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39127),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_335_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_hc_sig_LC_14_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_14_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_14_5_4  (
            .in0(N__36451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47982),
            .ce(),
            .sr(N__47273));
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_6_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_6_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_14_6_5  (
            .in0(N__36573),
            .in1(N__36553),
            .in2(N__47464),
            .in3(N__36441),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47974),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_14_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_14_8_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_14_8_1  (
            .in0(N__41205),
            .in1(N__34511),
            .in2(N__40729),
            .in3(N__40852),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47958),
            .ce(),
            .sr(N__47289));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_14_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_14_8_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_14_8_3  (
            .in0(N__40709),
            .in1(N__41447),
            .in2(N__35360),
            .in3(N__40850),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47958),
            .ce(),
            .sr(N__47289));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_14_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_14_8_5 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_14_8_5 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_14_8_5  (
            .in0(N__35252),
            .in1(N__42436),
            .in2(N__40728),
            .in3(N__40851),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47958),
            .ce(),
            .sr(N__47289));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_9_3  (
            .in0(N__41550),
            .in1(N__41442),
            .in2(N__41395),
            .in3(N__41488),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_11_LC_14_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_11_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_11_LC_14_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_11_LC_14_9_4  (
            .in0(N__41487),
            .in1(N__44284),
            .in2(N__41446),
            .in3(N__44305),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_5_LC_14_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_5_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_5_LC_14_9_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_5_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__41207),
            .in2(_gnd_net_),
            .in3(N__42475),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQI9C2_13_LC_14_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQI9C2_13_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQI9C2_13_LC_14_9_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQI9C2_13_LC_14_9_7  (
            .in0(N__41391),
            .in1(N__34187),
            .in2(N__34181),
            .in3(N__44227),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_14_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_14_10_0 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_14_10_0  (
            .in0(N__40666),
            .in1(N__44309),
            .in2(N__35095),
            .in3(N__40846),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47949),
            .ce(),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_14_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_14_10_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_14_10_1  (
            .in0(N__40847),
            .in1(N__44357),
            .in2(N__34606),
            .in3(N__40670),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47949),
            .ce(),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_14_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_14_10_5 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_14_10_5  (
            .in0(N__40848),
            .in1(N__34543),
            .in2(N__41711),
            .in3(N__40671),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47949),
            .ce(),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_14_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_14_10_6 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_14_10_6  (
            .in0(N__35488),
            .in1(N__41644),
            .in2(N__40716),
            .in3(N__40849),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47949),
            .ce(),
            .sr(N__47293));
    defparam \phase_controller_inst1.state_1_LC_14_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_14_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_14_11_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_1_LC_14_11_0  (
            .in0(N__34176),
            .in1(N__34379),
            .in2(N__34123),
            .in3(N__34346),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47939),
            .ce(),
            .sr(N__47299));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_14_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_14_11_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_14_11_2  (
            .in0(N__40653),
            .in1(N__34680),
            .in2(N__41555),
            .in3(N__40842),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47939),
            .ce(),
            .sr(N__47299));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_14_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_14_11_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_14_11_4  (
            .in0(N__40652),
            .in1(N__34486),
            .in2(_gnd_net_),
            .in3(N__40843),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47939),
            .ce(),
            .sr(N__47299));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_14_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_14_12_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_14_12_0  (
            .in0(N__37064),
            .in1(N__39659),
            .in2(N__39641),
            .in3(N__34472),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_12_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_12_1  (
            .in0(N__34259),
            .in1(N__38624),
            .in2(_gnd_net_),
            .in3(N__39221),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_1_LC_14_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_1_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_1_LC_14_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_1_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__34512),
            .in2(_gnd_net_),
            .in3(N__39759),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_14_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_14_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_14_12_3  (
            .in0(N__35090),
            .in1(N__34736),
            .in2(N__36746),
            .in3(N__34809),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_14_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_14_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_14_12_4  (
            .in0(N__34557),
            .in1(N__34672),
            .in2(N__35500),
            .in3(N__35089),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_12_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__34595),
            .in2(_gnd_net_),
            .in3(N__35304),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_14_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_14_12_6  (
            .in0(N__34808),
            .in1(N__35187),
            .in2(N__34741),
            .in3(N__35132),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_14_12_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__39677),
            .in2(_gnd_net_),
            .in3(N__34487),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__34451),
            .in2(_gnd_net_),
            .in3(N__34411),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_14_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_14_13_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_14_13_1  (
            .in0(N__40024),
            .in1(N__34463),
            .in2(N__34466),
            .in3(N__42908),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47922),
            .ce(),
            .sr(N__47313));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__34371),
            .in2(_gnd_net_),
            .in3(N__34340),
            .lcout(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_13_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_13_3  (
            .in0(N__34452),
            .in1(N__34345),
            .in2(N__34378),
            .in3(N__34412),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47922),
            .ce(),
            .sr(N__47313));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_13_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_13_4  (
            .in0(N__39957),
            .in1(N__40025),
            .in2(N__37358),
            .in3(N__40231),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47922),
            .ce(),
            .sr(N__47313));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_13_5 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_14_13_5  (
            .in0(N__34341),
            .in1(N__34314),
            .in2(N__34358),
            .in3(N__34293),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47922),
            .ce(),
            .sr(N__47313));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_14_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__39956),
            .in2(_gnd_net_),
            .in3(N__40230),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34298),
            .in3(N__34292),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_14_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_14_0  (
            .in0(N__39950),
            .in1(N__40239),
            .in2(N__40125),
            .in3(N__37331),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_14_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_14_1  (
            .in0(N__40233),
            .in1(N__40113),
            .in2(N__37310),
            .in3(N__39952),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_14_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_14_2  (
            .in0(N__39949),
            .in1(N__40238),
            .in2(N__40124),
            .in3(N__37085),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_14_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_14_3  (
            .in0(N__40234),
            .in1(N__40114),
            .in2(N__36998),
            .in3(N__39953),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_14_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_14_4  (
            .in0(N__39951),
            .in1(N__40240),
            .in2(N__40126),
            .in3(N__36953),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_14_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_14_5  (
            .in0(N__40236),
            .in1(N__40116),
            .in2(N__37193),
            .in3(N__39955),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_14_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_14_6  (
            .in0(N__39948),
            .in1(N__40237),
            .in2(N__40123),
            .in3(N__37109),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_14_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_14_7  (
            .in0(N__40235),
            .in1(N__40115),
            .in2(N__36863),
            .in3(N__39954),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47915),
            .ce(),
            .sr(N__47319));
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_14_15_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_0_LC_14_15_0  (
            .in0(N__34986),
            .in1(N__40463),
            .in2(N__35615),
            .in3(N__39592),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47911),
            .ce(N__39801),
            .sr(N__47325));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_15_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_15_1 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_14_15_1  (
            .in0(N__36417),
            .in1(N__35600),
            .in2(N__40531),
            .in3(N__34985),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47911),
            .ce(N__39801),
            .sr(N__47325));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_14_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_14_15_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_14_15_3  (
            .in0(N__40462),
            .in1(N__34903),
            .in2(_gnd_net_),
            .in3(N__34877),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_15_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_15_4 .LUT_INIT=16'b1000110011001100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_14_15_4  (
            .in0(N__39722),
            .in1(N__34843),
            .in2(N__34823),
            .in3(N__34771),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47911),
            .ce(N__39801),
            .sr(N__47325));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_14_15_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_14_15_6 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_14_15_6  (
            .in0(N__35598),
            .in1(N__40464),
            .in2(N__34820),
            .in3(N__34769),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47911),
            .ce(N__39801),
            .sr(N__47325));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_15_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_15_7 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_14_15_7  (
            .in0(N__34770),
            .in1(N__35599),
            .in2(N__40530),
            .in3(N__34737),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47911),
            .ce(N__39801),
            .sr(N__47325));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_14_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_14_16_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_14_16_0  (
            .in0(N__40475),
            .in1(N__34681),
            .in2(_gnd_net_),
            .in3(N__35009),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_14_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_14_16_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_14_16_1  (
            .in0(N__35010),
            .in1(N__40476),
            .in2(_gnd_net_),
            .in3(N__34649),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_14_16_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_14_16_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_14_16_2  (
            .in0(N__35584),
            .in1(N__34596),
            .in2(N__40534),
            .in3(N__35437),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_14_16_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_14_16_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_14_16_3  (
            .in0(N__35439),
            .in1(N__35586),
            .in2(N__34565),
            .in3(N__40486),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_14_16_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_14_16_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_14_16_4  (
            .in0(N__40478),
            .in1(N__35012),
            .in2(_gnd_net_),
            .in3(N__34513),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_16_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_16_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_14_16_5  (
            .in0(N__35011),
            .in1(N__40477),
            .in2(_gnd_net_),
            .in3(N__35364),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_14_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_14_16_6 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_14_16_6  (
            .in0(N__35583),
            .in1(N__35315),
            .in2(N__40533),
            .in3(N__35436),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_14_16_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_14_16_7 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_14_16_7  (
            .in0(N__35438),
            .in1(N__35585),
            .in2(N__35279),
            .in3(N__40485),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47905),
            .ce(N__39817),
            .sr(N__47337));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_17_0 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_14_17_0  (
            .in0(N__35221),
            .in1(N__40471),
            .in2(_gnd_net_),
            .in3(N__36799),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_14_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_14_17_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_14_17_2  (
            .in0(N__35451),
            .in1(N__35611),
            .in2(N__40537),
            .in3(N__35195),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_14_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_14_17_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_14_17_3  (
            .in0(N__35014),
            .in1(N__40497),
            .in2(_gnd_net_),
            .in3(N__35144),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_4  (
            .in0(N__40498),
            .in1(N__35015),
            .in2(_gnd_net_),
            .in3(N__39767),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_17_5 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_14_17_5  (
            .in0(N__35091),
            .in1(N__40502),
            .in2(N__35618),
            .in3(N__35452),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_17_6 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_17_6  (
            .in0(N__40496),
            .in1(N__35056),
            .in2(_gnd_net_),
            .in3(N__35013),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_14_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_14_17_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_14_17_7  (
            .in0(N__35610),
            .in1(N__35501),
            .in2(N__40532),
            .in3(N__35453),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47899),
            .ce(N__39818),
            .sr(N__47347));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__37649),
            .in2(N__37733),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__38381),
            .in2(_gnd_net_),
            .in3(N__35390),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__37685),
            .in2(N__38360),
            .in3(N__35387),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__38336),
            .in2(_gnd_net_),
            .in3(N__35384),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__38315),
            .in2(_gnd_net_),
            .in3(N__35381),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_18_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38294),
            .in3(N__35378),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__38269),
            .in2(_gnd_net_),
            .in3(N__35375),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__38239),
            .in2(_gnd_net_),
            .in3(N__35372),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__38218),
            .in2(_gnd_net_),
            .in3(N__35651),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__38548),
            .in2(_gnd_net_),
            .in3(N__35648),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__38527),
            .in2(_gnd_net_),
            .in3(N__35645),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__38506),
            .in2(_gnd_net_),
            .in3(N__35642),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__38485),
            .in2(_gnd_net_),
            .in3(N__35639),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__38464),
            .in2(_gnd_net_),
            .in3(N__35636),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__38443),
            .in2(_gnd_net_),
            .in3(N__35633),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_19_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38407),
            .in3(N__35624),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__38767),
            .in2(_gnd_net_),
            .in3(N__35621),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__38743),
            .in2(_gnd_net_),
            .in3(N__35711),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__38722),
            .in2(_gnd_net_),
            .in3(N__35708),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_14_21_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_14_21_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_14_21_0  (
            .in0(N__37842),
            .in1(N__38117),
            .in2(N__38012),
            .in3(N__35705),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_14_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_14_21_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_14_21_1  (
            .in0(N__38113),
            .in1(N__37991),
            .in2(N__37869),
            .in3(N__35699),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_14_21_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_14_21_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_14_21_2  (
            .in0(N__37843),
            .in1(N__38118),
            .in2(N__38013),
            .in3(N__35693),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_21_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_21_3  (
            .in0(N__38114),
            .in1(N__37992),
            .in2(N__37870),
            .in3(N__35687),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_21_4 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_21_4  (
            .in0(N__37844),
            .in1(N__35678),
            .in2(N__38014),
            .in3(N__38120),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_21_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_21_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_21_5  (
            .in0(N__38115),
            .in1(N__37993),
            .in2(N__37871),
            .in3(N__35669),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_21_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_21_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_21_6  (
            .in0(N__37845),
            .in1(N__38119),
            .in2(N__38015),
            .in3(N__35660),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_21_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_21_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_21_7  (
            .in0(N__38116),
            .in1(N__37994),
            .in2(N__37872),
            .in3(N__35759),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47879),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_14_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_14_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48334),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47871),
            .ce(N__43354),
            .sr(N__47384));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_14_22_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_14_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__43445),
            .in2(_gnd_net_),
            .in3(N__46823),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47871),
            .ce(N__43354),
            .sr(N__47384));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_23_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_23_0  (
            .in0(N__36316),
            .in1(N__36104),
            .in2(N__36055),
            .in3(N__35750),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47866),
            .ce(),
            .sr(N__47393));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_23_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_23_2  (
            .in0(N__36317),
            .in1(N__36105),
            .in2(N__36056),
            .in3(N__35744),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47866),
            .ce(),
            .sr(N__47393));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_23_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_23_3  (
            .in0(N__36103),
            .in1(N__36021),
            .in2(_gnd_net_),
            .in3(N__36315),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_14_23_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_14_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_14_23_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_14_23_5  (
            .in0(N__43585),
            .in1(N__43853),
            .in2(N__43732),
            .in3(N__37679),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47866),
            .ce(),
            .sr(N__47393));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_24_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_24_0  (
            .in0(N__36294),
            .in1(N__36155),
            .in2(N__36064),
            .in3(N__35735),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_24_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_24_1  (
            .in0(N__36034),
            .in1(N__36287),
            .in2(N__36181),
            .in3(N__35729),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_24_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_24_2  (
            .in0(N__36289),
            .in1(N__36144),
            .in2(N__36062),
            .in3(N__35723),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_24_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_24_3  (
            .in0(N__36035),
            .in1(N__36290),
            .in2(N__36182),
            .in3(N__35813),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_24_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_24_4  (
            .in0(N__36291),
            .in1(N__36148),
            .in2(N__36063),
            .in3(N__35807),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_24_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_24_5  (
            .in0(N__36036),
            .in1(N__36292),
            .in2(N__36183),
            .in3(N__35801),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_24_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_24_6  (
            .in0(N__36288),
            .in1(N__36143),
            .in2(N__36061),
            .in3(N__35795),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_24_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_24_7  (
            .in0(N__36037),
            .in1(N__36293),
            .in2(N__36184),
            .in3(N__35789),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47861),
            .ce(),
            .sr(N__47397));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_25_0 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_25_0  (
            .in0(N__36000),
            .in1(N__35783),
            .in2(N__36205),
            .in3(N__36318),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_25_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_25_1  (
            .in0(N__36322),
            .in1(N__36193),
            .in2(N__36052),
            .in3(N__35777),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_25_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_25_2  (
            .in0(N__36003),
            .in1(N__36325),
            .in2(N__36208),
            .in3(N__35771),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_25_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_25_3  (
            .in0(N__36324),
            .in1(N__36197),
            .in2(N__36053),
            .in3(N__35765),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_25_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_25_4  (
            .in0(N__36002),
            .in1(N__36323),
            .in2(N__36207),
            .in3(N__36350),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_25_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_25_5  (
            .in0(N__36321),
            .in1(N__36192),
            .in2(N__36051),
            .in3(N__36344),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_25_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_25_6  (
            .in0(N__36001),
            .in1(N__36319),
            .in2(N__36206),
            .in3(N__36338),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_25_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_25_7  (
            .in0(N__36320),
            .in1(N__36191),
            .in2(N__36050),
            .in3(N__36332),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47855),
            .ce(),
            .sr(N__47400));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_26_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_26_6 .LUT_INIT=16'b0100000001100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_26_6  (
            .in0(N__36326),
            .in1(N__36016),
            .in2(N__36209),
            .in3(N__39201),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47852),
            .ce(N__35861),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR1_LC_15_4_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_4_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_15_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35912),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47993),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_15_4_6.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_4_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_15_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35903),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47993),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_15_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_15_5_1 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_15_5_1  (
            .in0(N__36525),
            .in1(N__36507),
            .in2(_gnd_net_),
            .in3(N__36491),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__35879),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_tr_sig_LC_15_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_15_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36535),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(),
            .sr(N__47274));
    defparam \delay_measurement_inst.start_timer_hc_LC_15_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_6_5 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_15_6_5  (
            .in0(N__36575),
            .in1(N__36557),
            .in2(_gnd_net_),
            .in3(N__36440),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(),
            .sr(N__47274));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6  (
            .in0(N__39140),
            .in1(N__39126),
            .in2(_gnd_net_),
            .in3(N__39103),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(),
            .sr(N__47274));
    defparam \delay_measurement_inst.start_timer_tr_LC_15_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_6_7 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_15_6_7  (
            .in0(N__36534),
            .in1(N__36508),
            .in2(_gnd_net_),
            .in3(N__36489),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(),
            .sr(N__47274));
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_7_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_15_7_0  (
            .in0(N__36536),
            .in1(N__36512),
            .in2(N__47465),
            .in3(N__36490),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47975),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC1_LC_15_7_3.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_15_7_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_15_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_15_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36473),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47975),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_15_7_7.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_15_7_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_15_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_15_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36458),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47975),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_15_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_15_8_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_15_8_0 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_15_8_0  (
            .in0(N__40693),
            .in1(N__44078),
            .in2(N__36413),
            .in3(N__36704),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47966),
            .ce(),
            .sr(N__47286));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_8_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_8_1  (
            .in0(N__36645),
            .in1(N__36364),
            .in2(_gnd_net_),
            .in3(N__36596),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_338_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_15_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_15_8_2 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_15_8_2  (
            .in0(N__36597),
            .in1(N__36365),
            .in2(_gnd_net_),
            .in3(N__36646),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47966),
            .ce(),
            .sr(N__47286));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_9_0 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_9_0  (
            .in0(N__44355),
            .in1(N__44257),
            .in2(N__41554),
            .in3(N__42432),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITLCJ3_7_LC_15_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITLCJ3_7_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITLCJ3_7_LC_15_9_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITLCJ3_7_LC_15_9_1  (
            .in0(N__36629),
            .in1(N__41643),
            .in2(N__36650),
            .in3(N__41707),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__36647),
            .in2(_gnd_net_),
            .in3(N__36598),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_337_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_15_LC_15_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_15_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_15_LC_15_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_15_LC_15_9_6  (
            .in0(N__44080),
            .in1(N__44138),
            .in2(N__42010),
            .in3(N__44020),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_15_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_15_10_2 .LUT_INIT=16'b0101110100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_15_10_2  (
            .in0(N__42369),
            .in1(N__44081),
            .in2(N__36833),
            .in3(N__44149),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_13_LC_15_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_13_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_13_LC_15_10_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_13_LC_15_10_5  (
            .in0(N__36620),
            .in1(N__36614),
            .in2(N__39380),
            .in3(N__39365),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_15_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_15_10_6 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_15_10_6  (
            .in0(N__36608),
            .in1(N__42011),
            .in2(N__36602),
            .in3(N__43956),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36599),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB9F91_3_LC_15_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB9F91_3_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB9F91_3_LC_15_11_2 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB9F91_3_LC_15_11_2  (
            .in0(N__42470),
            .in1(N__42431),
            .in2(_gnd_net_),
            .in3(N__44014),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_c_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEB452_7_LC_15_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEB452_7_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEB452_7_LC_15_11_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEB452_7_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__41638),
            .in2(N__36851),
            .in3(N__41705),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH8A4_6_LC_15_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH8A4_6_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH8A4_6_LC_15_11_4 .LUT_INIT=16'b0010101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH8A4_6_LC_15_11_4  (
            .in0(N__44079),
            .in1(N__42391),
            .in2(N__36848),
            .in3(N__44015),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_7_LC_15_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_7_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_7_LC_15_11_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_7_LC_15_11_6  (
            .in0(N__41706),
            .in1(_gnd_net_),
            .in2(N__41645),
            .in3(N__44016),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_15_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_15_11_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_15_11_7  (
            .in0(N__41206),
            .in1(N__44356),
            .in2(_gnd_net_),
            .in3(N__41272),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_15_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_15_12_0  (
            .in0(N__36824),
            .in1(N__36762),
            .in2(N__36728),
            .in3(N__36741),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_15_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_15_12_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_15_12_1  (
            .in0(N__36763),
            .in1(N__40681),
            .in2(_gnd_net_),
            .in3(N__36696),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47940),
            .ce(),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_15_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_15_12_3 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_15_12_3  (
            .in0(N__36742),
            .in1(N__40684),
            .in2(N__44261),
            .in3(N__40792),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47940),
            .ce(),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_15_12_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_15_12_4  (
            .in0(N__40793),
            .in1(_gnd_net_),
            .in2(N__40721),
            .in3(N__36723),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47940),
            .ce(),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_15_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_15_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_15_12_5  (
            .in0(N__37076),
            .in1(N__40683),
            .in2(_gnd_net_),
            .in3(N__36697),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47940),
            .ce(),
            .sr(N__47300));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_15_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_15_12_6  (
            .in0(N__37075),
            .in1(N__39619),
            .in2(N__37058),
            .in3(N__39607),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_15_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_15_12_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_15_12_7  (
            .in0(N__37057),
            .in1(N__40682),
            .in2(_gnd_net_),
            .in3(N__40794),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47940),
            .ce(),
            .sr(N__47300));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__37043),
            .in2(N__37037),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__37010),
            .in2(_gnd_net_),
            .in3(N__36983),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__36980),
            .in2(N__36968),
            .in3(N__36947),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__36944),
            .in2(_gnd_net_),
            .in3(N__36911),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__36908),
            .in2(_gnd_net_),
            .in3(N__36878),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__36875),
            .in2(_gnd_net_),
            .in3(N__36854),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__37238),
            .in2(_gnd_net_),
            .in3(N__37208),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__37205),
            .in2(_gnd_net_),
            .in3(N__37184),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__37181),
            .in2(_gnd_net_),
            .in3(N__37157),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__40300),
            .in2(_gnd_net_),
            .in3(N__37154),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__37151),
            .in2(_gnd_net_),
            .in3(N__37124),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__37121),
            .in2(_gnd_net_),
            .in3(N__37103),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__40279),
            .in2(_gnd_net_),
            .in3(N__37100),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__37097),
            .in2(_gnd_net_),
            .in3(N__37079),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__40258),
            .in2(_gnd_net_),
            .in3(N__37376),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__37372),
            .in2(_gnd_net_),
            .in3(N__37349),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__37345),
            .in2(_gnd_net_),
            .in3(N__37325),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__37322),
            .in2(_gnd_net_),
            .in3(N__37301),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__39832),
            .in2(_gnd_net_),
            .in3(N__37298),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_16_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37295),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_16_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__37274),
            .in2(N__37286),
            .in3(N__45327),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_16_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__37259),
            .in2(N__37268),
            .in3(N__45295),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_16_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__37244),
            .in2(N__37253),
            .in3(N__45253),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_16_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__37481),
            .in2(N__37490),
            .in3(N__45220),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_16_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__37466),
            .in2(N__37475),
            .in3(N__45187),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_16_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__37451),
            .in2(N__37460),
            .in3(N__45151),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_16_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_16_7  (
            .in0(N__45643),
            .in1(N__37436),
            .in2(N__37445),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__37418),
            .in2(N__37430),
            .in3(N__45610),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__37400),
            .in2(N__37412),
            .in3(N__45581),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__37382),
            .in2(N__37394),
            .in3(N__45547),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_17_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__37628),
            .in2(N__37643),
            .in3(N__45518),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_17_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__37610),
            .in2(N__37622),
            .in3(N__45491),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_17_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__37592),
            .in2(N__37604),
            .in3(N__45464),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_17_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_17_6  (
            .in0(N__45889),
            .in1(N__37571),
            .in2(N__37586),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_17_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__37553),
            .in2(N__37565),
            .in3(N__45863),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__37532),
            .in2(N__37547),
            .in3(N__45836),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__37511),
            .in2(N__37526),
            .in3(N__45809),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__37496),
            .in2(N__37505),
            .in3(N__45782),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__37703),
            .in2(N__37697),
            .in3(N__45755),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37688),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_15_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_15_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__38191),
            .in2(_gnd_net_),
            .in3(N__38681),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_18_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_18_7  (
            .in0(N__43063),
            .in1(N__45328),
            .in2(_gnd_net_),
            .in3(N__43015),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_19_0 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_19_0  (
            .in0(N__37667),
            .in1(N__37841),
            .in2(N__38131),
            .in3(N__37938),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47893),
            .ce(),
            .sr(N__47355));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_19_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_19_1  (
            .in0(N__37840),
            .in1(N__38106),
            .in2(N__37978),
            .in3(N__37661),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47893),
            .ce(),
            .sr(N__47355));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_19_2 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_19_2  (
            .in0(N__37839),
            .in1(N__37934),
            .in2(N__38130),
            .in3(N__37655),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47893),
            .ce(),
            .sr(N__47355));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_15_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_15_19_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_15_19_3  (
            .in0(N__37933),
            .in1(N__37838),
            .in2(_gnd_net_),
            .in3(N__38105),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__38190),
            .in2(_gnd_net_),
            .in3(N__38680),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_20_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_20_0  (
            .in0(N__37858),
            .in1(N__38123),
            .in2(N__38009),
            .in3(N__38198),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_20_1  (
            .in0(N__38192),
            .in1(N__37729),
            .in2(_gnd_net_),
            .in3(N__38682),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_20_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_20_2  (
            .in0(N__37861),
            .in1(N__38007),
            .in2(N__38159),
            .in3(N__38129),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_15_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_15_20_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_15_20_3  (
            .in0(N__38156),
            .in1(N__37979),
            .in2(N__38132),
            .in3(N__37862),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_20_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_20_4  (
            .in0(N__37859),
            .in1(N__38124),
            .in2(N__38010),
            .in3(N__38150),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_20_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_20_5  (
            .in0(N__38121),
            .in1(N__37980),
            .in2(N__37873),
            .in3(N__38144),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_20_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_20_6  (
            .in0(N__37860),
            .in1(N__38125),
            .in2(N__38011),
            .in3(N__38138),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_20_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_20_7  (
            .in0(N__38122),
            .in1(N__37981),
            .in2(N__37874),
            .in3(N__37739),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47886),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_21_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__37709),
            .in2(N__40892),
            .in3(N__37725),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_21_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__38366),
            .in2(N__40910),
            .in3(N__38377),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_21_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__38342),
            .in2(N__41006),
            .in3(N__38353),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_21_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__38321),
            .in2(N__40862),
            .in3(N__38332),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_21_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__38300),
            .in2(N__40997),
            .in3(N__38311),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_21_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__38276),
            .in2(N__40883),
            .in3(N__38287),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_21_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__38255),
            .in2(N__40871),
            .in3(N__38270),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_21_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__38225),
            .in2(N__38249),
            .in3(N__38240),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_22_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__38204),
            .in2(N__40937),
            .in3(N__38219),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_22_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_22_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_22_1  (
            .in0(N__38549),
            .in1(N__38534),
            .in2(N__40985),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_22_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__38513),
            .in2(N__40973),
            .in3(N__38528),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_22_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__38492),
            .in2(N__40949),
            .in3(N__38507),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_22_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_22_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_22_4  (
            .in0(N__38486),
            .in1(N__38471),
            .in2(N__40958),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_22_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__38450),
            .in2(N__43373),
            .in3(N__38465),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_22_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_22_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_22_6  (
            .in0(N__38444),
            .in1(N__40898),
            .in2(N__38429),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_22_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__38387),
            .in2(N__38420),
            .in3(N__38408),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_23_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__38753),
            .in2(N__38642),
            .in3(N__38771),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_23_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__38729),
            .in2(N__38633),
            .in3(N__38747),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_23_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_23_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_23_2  (
            .in0(N__38723),
            .in1(N__38708),
            .in2(N__40928),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_23_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38702),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_15_23_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_15_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48373),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47872),
            .ce(N__43353),
            .sr(N__47385));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_15_23_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_15_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48409),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47872),
            .ce(N__43353),
            .sr(N__47385));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__38597),
            .in2(N__41114),
            .in3(N__38613),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__40919),
            .in2(N__38579),
            .in3(N__38590),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__38555),
            .in2(N__41129),
            .in3(N__38566),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__38897),
            .in2(N__41141),
            .in3(N__38908),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_24_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_24_4  (
            .in0(N__38890),
            .in1(N__38879),
            .in2(N__41036),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__41147),
            .in2(N__38861),
            .in3(N__38872),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_24_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_24_6  (
            .in0(N__38851),
            .in1(N__38840),
            .in2(N__41105),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_24_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_24_7  (
            .in0(N__38833),
            .in1(N__38822),
            .in2(N__41045),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__38795),
            .in2(N__41339),
            .in3(N__38812),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_25_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_25_1  (
            .in0(N__38788),
            .in1(N__38777),
            .in2(N__41057),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__39062),
            .in2(N__41090),
            .in3(N__39073),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_25_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_25_3  (
            .in0(N__39055),
            .in1(N__39044),
            .in2(N__41288),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_25_4  (
            .in0(_gnd_net_),
            .in1(N__39026),
            .in2(N__41330),
            .in3(N__39037),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(N__39008),
            .in2(N__41321),
            .in3(N__39019),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__43136),
            .in2(N__38990),
            .in3(N__39001),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_25_7  (
            .in0(_gnd_net_),
            .in1(N__38951),
            .in2(N__38981),
            .in3(N__38969),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__38933),
            .in2(N__39167),
            .in3(N__38944),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__38915),
            .in2(N__39158),
            .in3(N__38926),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_26_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__39230),
            .in2(N__39149),
            .in3(N__39241),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_26_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39224),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_26_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_26_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48377),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47856),
            .ce(N__43103),
            .sr(N__47401));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_26_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_26_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_15_26_5  (
            .in0(N__48410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47856),
            .ce(N__43103),
            .sr(N__47401));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_26_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48059),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47856),
            .ce(N__43103),
            .sr(N__47401));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_6_2 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_6_2  (
            .in0(N__39102),
            .in1(N__39139),
            .in2(_gnd_net_),
            .in3(N__39128),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_336_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39101),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0  (
            .in0(N__39548),
            .in1(N__41247),
            .in2(_gnd_net_),
            .in3(N__39080),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1  (
            .in0(N__39504),
            .in1(N__44373),
            .in2(_gnd_net_),
            .in3(N__39077),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2  (
            .in0(N__39549),
            .in1(N__41226),
            .in2(_gnd_net_),
            .in3(N__39269),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3  (
            .in0(N__39505),
            .in1(N__41169),
            .in2(_gnd_net_),
            .in3(N__39266),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4  (
            .in0(N__39550),
            .in1(N__41730),
            .in2(_gnd_net_),
            .in3(N__39263),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5  (
            .in0(N__39506),
            .in1(N__41664),
            .in2(_gnd_net_),
            .in3(N__39260),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6  (
            .in0(N__39551),
            .in1(N__41598),
            .in2(_gnd_net_),
            .in3(N__39257),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7  (
            .in0(N__39507),
            .in1(N__41574),
            .in2(_gnd_net_),
            .in3(N__39254),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__47984),
            .ce(N__39405),
            .sr(N__47275));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0  (
            .in0(N__39539),
            .in1(N__41514),
            .in2(_gnd_net_),
            .in3(N__39251),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1  (
            .in0(N__39517),
            .in1(N__41466),
            .in2(_gnd_net_),
            .in3(N__39248),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2  (
            .in0(N__39536),
            .in1(N__41415),
            .in2(_gnd_net_),
            .in3(N__39245),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3  (
            .in0(N__39514),
            .in1(N__41361),
            .in2(_gnd_net_),
            .in3(N__39296),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4  (
            .in0(N__39537),
            .in1(N__42045),
            .in2(_gnd_net_),
            .in3(N__39293),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5  (
            .in0(N__39515),
            .in1(N__41958),
            .in2(_gnd_net_),
            .in3(N__39290),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6  (
            .in0(N__39538),
            .in1(N__41934),
            .in2(_gnd_net_),
            .in3(N__39287),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7  (
            .in0(N__39516),
            .in1(N__41910),
            .in2(_gnd_net_),
            .in3(N__39284),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__47976),
            .ce(N__39423),
            .sr(N__47278));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0  (
            .in0(N__39544),
            .in1(N__41886),
            .in2(_gnd_net_),
            .in3(N__39281),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1  (
            .in0(N__39540),
            .in1(N__41862),
            .in2(_gnd_net_),
            .in3(N__39278),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2  (
            .in0(N__39545),
            .in1(N__41820),
            .in2(_gnd_net_),
            .in3(N__39275),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3  (
            .in0(N__39541),
            .in1(N__41775),
            .in2(_gnd_net_),
            .in3(N__39272),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4  (
            .in0(N__39546),
            .in1(N__42318),
            .in2(_gnd_net_),
            .in3(N__39323),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5  (
            .in0(N__39542),
            .in1(N__42288),
            .in2(_gnd_net_),
            .in3(N__39320),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6  (
            .in0(N__39547),
            .in1(N__42258),
            .in2(_gnd_net_),
            .in3(N__39317),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7  (
            .in0(N__39543),
            .in1(N__42228),
            .in2(_gnd_net_),
            .in3(N__39314),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__47967),
            .ce(N__39425),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0  (
            .in0(N__39508),
            .in1(N__42198),
            .in2(_gnd_net_),
            .in3(N__39311),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__47959),
            .ce(N__39424),
            .sr(N__47290));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1  (
            .in0(N__39512),
            .in1(N__42168),
            .in2(_gnd_net_),
            .in3(N__39308),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__47959),
            .ce(N__39424),
            .sr(N__47290));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2  (
            .in0(N__39509),
            .in1(N__42138),
            .in2(_gnd_net_),
            .in3(N__39305),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__47959),
            .ce(N__39424),
            .sr(N__47290));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3  (
            .in0(N__39513),
            .in1(N__42093),
            .in2(_gnd_net_),
            .in3(N__39302),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__47959),
            .ce(N__39424),
            .sr(N__47290));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4  (
            .in0(N__39510),
            .in1(N__42118),
            .in2(_gnd_net_),
            .in3(N__39299),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__47959),
            .ce(N__39424),
            .sr(N__47290));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5  (
            .in0(N__42073),
            .in1(N__39511),
            .in2(_gnd_net_),
            .in3(N__39428),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47959),
            .ce(N__39424),
            .sr(N__47290));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVU8G_23_LC_16_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVU8G_23_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVU8G_23_LC_16_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVU8G_23_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__42269),
            .in2(_gnd_net_),
            .in3(N__42299),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_25_LC_16_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_25_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_25_LC_16_11_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_25_LC_16_11_1  (
            .in0(N__42209),
            .in1(N__42239),
            .in2(N__39389),
            .in3(N__39371),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII0UL_14_LC_16_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII0UL_14_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII0UL_14_LC_16_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII0UL_14_LC_16_11_3  (
            .in0(N__44071),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44134),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHOP1_7_LC_16_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHOP1_7_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHOP1_7_LC_16_11_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHOP1_7_LC_16_11_4  (
            .in0(N__41698),
            .in1(N__41642),
            .in2(N__39386),
            .in3(N__44182),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRLFA3_15_LC_16_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRLFA3_15_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRLFA3_15_LC_16_11_5 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRLFA3_15_LC_16_11_5  (
            .in0(N__44184),
            .in1(N__42012),
            .in2(N__39383),
            .in3(N__43950),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_16_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_16_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_16_11_6  (
            .in0(N__41797),
            .in1(N__41836),
            .in2(N__41752),
            .in3(N__44183),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_11_7  (
            .in0(N__42104),
            .in1(N__42149),
            .in2(N__42059),
            .in3(N__42179),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_12_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_12_4  (
            .in0(N__39364),
            .in1(N__41756),
            .in2(N__41843),
            .in3(N__41801),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto30_2 ),
            .ltout(\delay_measurement_inst.delay_hc_reg3lto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVBSED_31_LC_16_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVBSED_31_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVBSED_31_LC_16_12_5 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVBSED_31_LC_16_12_5  (
            .in0(N__39779),
            .in1(N__44185),
            .in2(N__39773),
            .in3(N__42344),
            .lcout(\delay_measurement_inst.delay_hc_reg3 ),
            .ltout(\delay_measurement_inst.delay_hc_reg3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_16_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_16_12_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_16_12_6  (
            .in0(N__40702),
            .in1(N__42474),
            .in2(N__39770),
            .in3(N__39758),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47950),
            .ce(),
            .sr(N__47294));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_16_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_16_13_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_16_13_0 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_16_13_0  (
            .in0(N__40697),
            .in1(N__44145),
            .in2(N__39712),
            .in3(N__40785),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_16_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_16_13_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_16_13_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_16_13_1  (
            .in0(N__40786),
            .in1(N__40698),
            .in2(_gnd_net_),
            .in3(N__39673),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_16_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_16_13_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_16_13_2  (
            .in0(N__40695),
            .in1(N__39655),
            .in2(_gnd_net_),
            .in3(N__40787),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_16_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_16_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_16_13_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_16_13_3  (
            .in0(N__40788),
            .in1(N__40699),
            .in2(_gnd_net_),
            .in3(N__39634),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_16_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_16_13_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_16_13_4  (
            .in0(N__40696),
            .in1(N__39620),
            .in2(_gnd_net_),
            .in3(N__40789),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_16_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_16_13_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_16_13_5  (
            .in0(N__40790),
            .in1(N__40700),
            .in2(_gnd_net_),
            .in3(N__39608),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_16_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_16_13_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_16_13_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_16_13_6  (
            .in0(N__40694),
            .in1(N__39581),
            .in2(_gnd_net_),
            .in3(N__40784),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_16_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_16_13_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_16_13_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_16_13_7  (
            .in0(N__40791),
            .in1(N__40701),
            .in2(_gnd_net_),
            .in3(N__40358),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47941),
            .ce(),
            .sr(N__47301));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_16_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_16_14_0 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_16_14_0  (
            .in0(N__39962),
            .in1(N__40307),
            .in2(N__40120),
            .in3(N__40244),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47930),
            .ce(),
            .sr(N__47307));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_16_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_16_14_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_16_14_2  (
            .in0(N__39963),
            .in1(N__40242),
            .in2(N__40121),
            .in3(N__40286),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47930),
            .ce(),
            .sr(N__47307));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_16_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_16_14_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_16_14_6  (
            .in0(N__39964),
            .in1(N__40243),
            .in2(N__40122),
            .in3(N__40265),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47930),
            .ce(),
            .sr(N__47307));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_16_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_16_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_16_14_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_16_14_7  (
            .in0(N__40241),
            .in1(N__40090),
            .in2(N__39974),
            .in3(N__39965),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47930),
            .ce(),
            .sr(N__47307));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_16_15_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_16_15_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_16_15_3  (
            .in0(N__43714),
            .in1(N__43583),
            .in2(_gnd_net_),
            .in3(N__43852),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_16_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_16_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_16_16_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_16_16_1  (
            .in0(N__43854),
            .in1(N__43584),
            .in2(N__43724),
            .in3(N__45632),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47916),
            .ce(),
            .sr(N__47320));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_16_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_16_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_16_17_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_16_17_0  (
            .in0(N__43823),
            .in1(N__43558),
            .in2(N__43721),
            .in3(N__45284),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_16_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_16_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_16_17_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_16_17_1  (
            .in0(N__43556),
            .in1(N__43703),
            .in2(N__45599),
            .in3(N__43829),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_16_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_16_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_16_17_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_16_17_2  (
            .in0(N__43824),
            .in1(N__43559),
            .in2(N__43722),
            .in3(N__45242),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_16_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_16_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_16_17_3 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_16_17_3  (
            .in0(N__43554),
            .in1(N__43701),
            .in2(N__45176),
            .in3(N__43827),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_16_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_16_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_16_17_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_16_17_4  (
            .in0(N__43822),
            .in1(N__43557),
            .in2(N__43720),
            .in3(N__45878),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_16_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_16_17_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_16_17_5  (
            .in0(N__43555),
            .in1(N__43702),
            .in2(N__45668),
            .in3(N__43828),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_16_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_16_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_16_17_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_16_17_6  (
            .in0(N__43825),
            .in1(N__43560),
            .in2(N__43723),
            .in3(N__45209),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_16_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_16_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_16_17_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_16_17_7  (
            .in0(N__43553),
            .in1(N__43700),
            .in2(N__45536),
            .in3(N__43826),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47912),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_16_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_16_18_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__43564),
            .in2(_gnd_net_),
            .in3(N__43834),
            .lcout(\phase_controller_slave.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_16_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_16_18_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_16_18_4  (
            .in0(N__43835),
            .in1(_gnd_net_),
            .in2(N__43586),
            .in3(N__43660),
            .lcout(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_19_3 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_19_3  (
            .in0(N__48260),
            .in1(N__48505),
            .in2(_gnd_net_),
            .in3(N__45950),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47900),
            .ce(N__47518),
            .sr(N__47348));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_19_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_19_6  (
            .in0(N__48506),
            .in1(N__48261),
            .in2(_gnd_net_),
            .in3(N__45968),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47900),
            .ce(N__47518),
            .sr(N__47348));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_16_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_16_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_16_20_0  (
            .in0(N__41304),
            .in1(N__48459),
            .in2(N__46678),
            .in3(N__41073),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_16_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_16_20_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40913),
            .in3(N__41019),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_20_5 .LUT_INIT=16'b0101010100000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_20_5  (
            .in0(N__42932),
            .in1(N__48504),
            .in2(N__48281),
            .in3(N__46034),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47894),
            .ce(N__47519),
            .sr(N__47356));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_16_21_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_16_21_0 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_16_21_0  (
            .in0(N__43244),
            .in1(N__43186),
            .in2(N__46432),
            .in3(N__43407),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_16_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_16_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__45712),
            .in2(_gnd_net_),
            .in3(N__46182),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_16_21_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_16_21_2 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_16_21_2  (
            .in0(N__43243),
            .in1(N__43185),
            .in2(N__46060),
            .in3(N__43406),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_16_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_16_21_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_6_LC_16_21_3  (
            .in0(N__43411),
            .in1(N__46615),
            .in2(_gnd_net_),
            .in3(N__43190),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_16_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_16_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__46759),
            .in2(_gnd_net_),
            .in3(N__43412),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_16_21_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_16_21_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_16_21_5  (
            .in0(N__43409),
            .in1(N__43188),
            .in2(_gnd_net_),
            .in3(N__46564),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_16_21_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_16_21_6 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_16_21_6  (
            .in0(N__43187),
            .in1(N__43408),
            .in2(N__46888),
            .in3(N__43263),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_16_21_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_16_21_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_16_21_7  (
            .in0(N__43410),
            .in1(N__43189),
            .in2(_gnd_net_),
            .in3(N__46945),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47887),
            .ce(N__43352),
            .sr(N__47365));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_16_22_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_16_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__43299),
            .in2(_gnd_net_),
            .in3(N__41080),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47883),
            .ce(N__43348),
            .sr(N__47374));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_16_22_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_16_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_16_22_1  (
            .in0(N__43300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48466),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47883),
            .ce(N__43348),
            .sr(N__47374));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_16_22_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_16_22_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_16_22_3  (
            .in0(N__43302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46674),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47883),
            .ce(N__43348),
            .sr(N__47374));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_16_22_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_16_22_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_16_22_4  (
            .in0(N__41311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43301),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47883),
            .ce(N__43348),
            .sr(N__47374));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_16_22_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_16_22_6 .LUT_INIT=16'b1101110011011101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_16_22_6  (
            .in0(N__43303),
            .in1(N__41027),
            .in2(N__46184),
            .in3(N__43218),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47883),
            .ce(N__43348),
            .sr(N__47374));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_22_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48054),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47883),
            .ce(N__43348),
            .sr(N__47374));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_23_0 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_16_23_0  (
            .in0(N__43161),
            .in1(N__43435),
            .in2(N__46433),
            .in3(N__43237),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47880),
            .ce(N__43094),
            .sr(N__47380));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_23_1 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_16_23_1  (
            .in0(N__43438),
            .in1(N__43164),
            .in2(_gnd_net_),
            .in3(N__46619),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47880),
            .ce(N__43094),
            .sr(N__47380));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_23_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_16_23_2  (
            .in0(N__43163),
            .in1(N__46568),
            .in2(_gnd_net_),
            .in3(N__43437),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47880),
            .ce(N__43094),
            .sr(N__47380));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_23_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_16_23_3  (
            .in0(N__43436),
            .in1(N__43162),
            .in2(N__46889),
            .in3(N__43265),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47880),
            .ce(N__43094),
            .sr(N__47380));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_23_6 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_16_23_6  (
            .in0(N__43160),
            .in1(N__43434),
            .in2(N__46067),
            .in3(N__43236),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47880),
            .ce(N__43094),
            .sr(N__47380));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_16_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_16_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(N__43440),
            .in2(_gnd_net_),
            .in3(N__46763),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(N__43110),
            .sr(N__47386));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_24_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_16_24_1  (
            .in0(N__43297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48467),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(N__43110),
            .sr(N__47386));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(N__43296),
            .in2(_gnd_net_),
            .in3(N__41081),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(N__43110),
            .sr(N__47386));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_24_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_16_24_3  (
            .in0(N__43441),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46822),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(N__43110),
            .sr(N__47386));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_24_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_16_24_6  (
            .in0(N__43165),
            .in1(N__46946),
            .in2(_gnd_net_),
            .in3(N__43439),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(N__43110),
            .sr(N__47386));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_24_7 .LUT_INIT=16'b1111111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_16_24_7  (
            .in0(N__43298),
            .in1(N__46183),
            .in2(N__43223),
            .in3(N__41026),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(N__43110),
            .sr(N__47386));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_25_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_16_25_2  (
            .in0(N__43310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46679),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__43123),
            .sr(N__47394));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_25_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_16_25_3  (
            .in0(N__45713),
            .in1(N__46181),
            .in2(_gnd_net_),
            .in3(N__46318),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__43123),
            .sr(N__47394));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_25_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__43309),
            .in2(_gnd_net_),
            .in3(N__41312),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__43123),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__41249),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47991),
            .ce(N__44328),
            .sr(N__47272));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__41248),
            .in2(N__41228),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__44374),
            .in2(N__41171),
            .in3(N__41231),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__41227),
            .in2(N__41732),
            .in3(N__41174),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__41170),
            .in2(N__41666),
            .in3(N__41150),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__41731),
            .in2(N__41600),
            .in3(N__41669),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__41665),
            .in2(N__41576),
            .in3(N__41603),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__41599),
            .in2(N__41516),
            .in3(N__41579),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__41575),
            .in2(N__41468),
            .in3(N__41519),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47985),
            .ce(N__44329),
            .sr(N__47276));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__41515),
            .in2(N__41417),
            .in3(N__41471),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__41467),
            .in2(N__41363),
            .in3(N__41420),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__41416),
            .in2(N__42047),
            .in3(N__41366),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__41362),
            .in2(N__41960),
            .in3(N__41342),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__42046),
            .in2(N__41936),
            .in3(N__41963),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__41959),
            .in2(N__41912),
            .in3(N__41939),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__41935),
            .in2(N__41888),
            .in3(N__41915),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__41911),
            .in2(N__41864),
            .in3(N__41891),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47977),
            .ce(N__44330),
            .sr(N__47279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__41887),
            .in2(N__41822),
            .in3(N__41867),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__41863),
            .in2(N__41777),
            .in3(N__41825),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__41821),
            .in2(N__42320),
            .in3(N__41780),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__41776),
            .in2(N__42290),
            .in3(N__41735),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__42319),
            .in2(N__42260),
            .in3(N__42293),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__42289),
            .in2(N__42230),
            .in3(N__42263),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__42259),
            .in2(N__42200),
            .in3(N__42233),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__42229),
            .in2(N__42170),
            .in3(N__42203),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47968),
            .ce(N__44331),
            .sr(N__47288));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__42199),
            .in2(N__42140),
            .in3(N__42173),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47960),
            .ce(N__44333),
            .sr(N__47291));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__42169),
            .in2(N__42095),
            .in3(N__42143),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47960),
            .ce(N__44333),
            .sr(N__47291));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__42139),
            .in2(N__42119),
            .in3(N__42098),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47960),
            .ce(N__44333),
            .sr(N__47291));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__42094),
            .in2(N__42074),
            .in3(N__42050),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47960),
            .ce(N__44333),
            .sr(N__47291));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42479),
            .lcout(\delay_measurement_inst.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47960),
            .ce(N__44333),
            .sr(N__47291));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4_3_LC_17_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4_3_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4_3_LC_17_12_2 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4_3_LC_17_12_2  (
            .in0(N__42476),
            .in1(N__42437),
            .in2(N__42401),
            .in3(N__43907),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4KK27_3_LC_17_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4KK27_3_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4KK27_3_LC_17_12_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4KK27_3_LC_17_12_3  (
            .in0(N__44090),
            .in1(N__42379),
            .in2(N__42347),
            .in3(N__43943),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_13_0  (
            .in0(N__42717),
            .in1(N__43896),
            .in2(_gnd_net_),
            .in3(N__42338),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_13_1  (
            .in0(N__42733),
            .in1(N__43875),
            .in2(_gnd_net_),
            .in3(N__42335),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_13_2  (
            .in0(N__42718),
            .in1(N__44619),
            .in2(_gnd_net_),
            .in3(N__42332),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_13_3  (
            .in0(N__42734),
            .in1(N__44592),
            .in2(_gnd_net_),
            .in3(N__42329),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_13_4  (
            .in0(N__42719),
            .in1(N__44566),
            .in2(_gnd_net_),
            .in3(N__42326),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_13_5  (
            .in0(N__42735),
            .in1(N__44542),
            .in2(_gnd_net_),
            .in3(N__42323),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_13_6  (
            .in0(N__42716),
            .in1(N__44514),
            .in2(_gnd_net_),
            .in3(N__42506),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_13_7  (
            .in0(N__42736),
            .in1(N__44482),
            .in2(_gnd_net_),
            .in3(N__42503),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__47951),
            .ce(N__42590),
            .sr(N__47295));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_14_0  (
            .in0(N__42711),
            .in1(N__44457),
            .in2(_gnd_net_),
            .in3(N__42500),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_14_1  (
            .in0(N__42723),
            .in1(N__44431),
            .in2(_gnd_net_),
            .in3(N__42497),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_14_2  (
            .in0(N__42708),
            .in1(N__44400),
            .in2(_gnd_net_),
            .in3(N__42494),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_14_3  (
            .in0(N__42720),
            .in1(N__44835),
            .in2(_gnd_net_),
            .in3(N__42491),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_14_4  (
            .in0(N__42709),
            .in1(N__44808),
            .in2(_gnd_net_),
            .in3(N__42488),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_14_5  (
            .in0(N__42721),
            .in1(N__44781),
            .in2(_gnd_net_),
            .in3(N__42485),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_14_6  (
            .in0(N__42710),
            .in1(N__44760),
            .in2(_gnd_net_),
            .in3(N__42482),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_14_7  (
            .in0(N__42722),
            .in1(N__44739),
            .in2(_gnd_net_),
            .in3(N__42533),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__47942),
            .ce(N__42591),
            .sr(N__47302));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_15_0  (
            .in0(N__42712),
            .in1(N__44715),
            .in2(_gnd_net_),
            .in3(N__42530),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_15_1  (
            .in0(N__42737),
            .in1(N__44688),
            .in2(_gnd_net_),
            .in3(N__42527),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_15_2  (
            .in0(N__42713),
            .in1(N__44652),
            .in2(_gnd_net_),
            .in3(N__42524),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_15_3  (
            .in0(N__42738),
            .in1(N__45132),
            .in2(_gnd_net_),
            .in3(N__42521),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_15_4  (
            .in0(N__42714),
            .in1(N__45100),
            .in2(_gnd_net_),
            .in3(N__42518),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_15_5  (
            .in0(N__42739),
            .in1(N__45066),
            .in2(_gnd_net_),
            .in3(N__42515),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_15_6  (
            .in0(N__42715),
            .in1(N__45027),
            .in2(_gnd_net_),
            .in3(N__42512),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_15_7  (
            .in0(N__42740),
            .in1(N__45000),
            .in2(_gnd_net_),
            .in3(N__42509),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__47931),
            .ce(N__42599),
            .sr(N__47308));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_16_0  (
            .in0(N__42702),
            .in1(N__44967),
            .in2(_gnd_net_),
            .in3(N__42755),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__47923),
            .ce(N__42595),
            .sr(N__47314));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_16_1  (
            .in0(N__42706),
            .in1(N__44931),
            .in2(_gnd_net_),
            .in3(N__42752),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__47923),
            .ce(N__42595),
            .sr(N__47314));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_16_2  (
            .in0(N__42703),
            .in1(N__44871),
            .in2(_gnd_net_),
            .in3(N__42749),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__47923),
            .ce(N__42595),
            .sr(N__47314));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_16_3  (
            .in0(N__42707),
            .in1(N__45435),
            .in2(_gnd_net_),
            .in3(N__42746),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__47923),
            .ce(N__42595),
            .sr(N__47314));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_16_4  (
            .in0(N__42704),
            .in1(N__44893),
            .in2(_gnd_net_),
            .in3(N__42743),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__47923),
            .ce(N__42595),
            .sr(N__47314));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_16_5  (
            .in0(N__45415),
            .in1(N__42705),
            .in2(_gnd_net_),
            .in3(N__42602),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47923),
            .ce(N__42595),
            .sr(N__47314));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_17_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_17_17_0 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_17_17_0  (
            .in0(N__46348),
            .in1(N__46028),
            .in2(_gnd_net_),
            .in3(N__45925),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_17_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_17_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_17_17_1  (
            .in0(N__44948),
            .in1(N__44984),
            .in2(N__44909),
            .in3(N__45011),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_17_5  (
            .in0(N__45086),
            .in1(N__45116),
            .in2(N__45050),
            .in3(N__44636),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_17_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_17_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_17_17_6  (
            .in0(N__44669),
            .in1(N__42956),
            .in2(N__42950),
            .in3(N__42938),
            .lcout(\delay_measurement_inst.N_358 ),
            .ltout(\delay_measurement_inst.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_17_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_17_17_7 .LUT_INIT=16'b0000111100000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_17_17_7  (
            .in0(N__46277),
            .in1(N__42947),
            .in2(N__42941),
            .in3(N__46213),
            .lcout(\delay_measurement_inst.N_324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_17_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_17_18_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__45401),
            .in2(_gnd_net_),
            .in3(N__44855),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_18_1  (
            .in0(N__43061),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43022),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_17_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_17_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_17_18_3  (
            .in0(N__43062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43023),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_17_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_17_18_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_17_18_5  (
            .in0(N__46029),
            .in1(N__45926),
            .in2(N__46276),
            .in3(N__48080),
            .lcout(\delay_measurement_inst.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_17_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_17_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__42823),
            .in2(_gnd_net_),
            .in3(N__42862),
            .lcout(),
            .ltout(\phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_LC_17_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_17_19_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_17_19_1  (
            .in0(N__43664),
            .in1(N__42923),
            .in2(N__42911),
            .in3(N__42903),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47906),
            .ce(),
            .sr(N__47338));
    defparam \phase_controller_slave.state_2_LC_17_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_17_19_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_slave.state_2_LC_17_19_3  (
            .in0(N__42863),
            .in1(N__42774),
            .in2(N__42827),
            .in3(N__42980),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47906),
            .ce(),
            .sr(N__47338));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_19_4 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_19_4  (
            .in0(N__43568),
            .in1(N__43665),
            .in2(N__43856),
            .in3(N__45500),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47906),
            .ce(),
            .sr(N__47338));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_17_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_17_19_5 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_17_19_5  (
            .in0(N__42981),
            .in1(N__43064),
            .in2(N__43043),
            .in3(N__43034),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47906),
            .ce(),
            .sr(N__47338));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_20_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_20_0  (
            .in0(N__43569),
            .in1(N__43842),
            .in2(N__43710),
            .in3(N__45473),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_20_1 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_20_1  (
            .in0(N__45563),
            .in1(N__43573),
            .in2(N__43855),
            .in3(N__43681),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_20_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_20_2  (
            .in0(N__43571),
            .in1(N__43844),
            .in2(N__43712),
            .in3(N__45845),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_20_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_20_3  (
            .in0(N__43839),
            .in1(N__43666),
            .in2(N__43587),
            .in3(N__45818),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_20_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_20_4  (
            .in0(N__43570),
            .in1(N__43843),
            .in2(N__43711),
            .in3(N__45446),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_20_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_20_5  (
            .in0(N__43840),
            .in1(N__43667),
            .in2(N__43588),
            .in3(N__45791),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_20_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_20_6  (
            .in0(N__43572),
            .in1(N__43845),
            .in2(N__43713),
            .in3(N__45764),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_20_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_20_7  (
            .in0(N__43841),
            .in1(N__43668),
            .in2(N__43589),
            .in3(N__45734),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47901),
            .ce(),
            .sr(N__47349));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_17_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_17_21_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_17_21_2  (
            .in0(N__46312),
            .in1(N__46941),
            .in2(N__46177),
            .in3(N__46563),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_17_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_17_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_17_21_3  (
            .in0(N__48299),
            .in1(N__45724),
            .in2(N__43463),
            .in3(N__43456),
            .lcout(\phase_controller_inst1.stoper_tr.N_279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_17_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_17_21_7 .LUT_INIT=16'b1011101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_17_21_7  (
            .in0(N__45693),
            .in1(N__46155),
            .in2(N__43460),
            .in3(N__46313),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_17_22_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_17_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_17_22_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_17_22_3  (
            .in0(N__45695),
            .in1(N__46173),
            .in2(_gnd_net_),
            .in3(N__46317),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47888),
            .ce(N__43358),
            .sr(N__47366));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_17_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_17_23_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_17_23_3  (
            .in0(N__45694),
            .in1(N__46179),
            .in2(_gnd_net_),
            .in3(N__46319),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_17_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_17_23_6 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_17_23_6  (
            .in0(N__46884),
            .in1(N__46422),
            .in2(_gnd_net_),
            .in3(N__43264),
            .lcout(\phase_controller_inst1.stoper_tr.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_17_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_17_23_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_17_23_7  (
            .in0(N__45728),
            .in1(N__43222),
            .in2(_gnd_net_),
            .in3(N__46178),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(N__45708),
            .in2(_gnd_net_),
            .in3(N__46180),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47874),
            .ce(N__43124),
            .sr(N__47387));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44381),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47986),
            .ce(N__44332),
            .sr(N__47277));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_18_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_18_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_18_10_1  (
            .in0(N__44298),
            .in1(N__44277),
            .in2(N__44250),
            .in3(N__44220),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITS8G_14_LC_18_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITS8G_14_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITS8G_14_LC_18_11_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITS8G_14_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__44181),
            .in2(_gnd_net_),
            .in3(N__44133),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA5CC2_6_LC_18_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA5CC2_6_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA5CC2_6_LC_18_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA5CC2_6_LC_18_11_7  (
            .in0(N__44067),
            .in1(N__44013),
            .in2(N__43970),
            .in3(N__43928),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43900),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47952),
            .ce(N__45373),
            .sr(N__47296));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43879),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47952),
            .ce(N__45373),
            .sr(N__47296));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__43901),
            .in2(N__44626),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__43880),
            .in2(N__44599),
            .in3(N__43859),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__44572),
            .in2(N__44627),
            .in3(N__44603),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__44548),
            .in2(N__44600),
            .in3(N__44576),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__44573),
            .in2(N__44525),
            .in3(N__44552),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__44549),
            .in2(N__44494),
            .in3(N__44528),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__44524),
            .in2(N__44461),
            .in3(N__44498),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__44430),
            .in2(N__44495),
            .in3(N__44468),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47943),
            .ce(N__45389),
            .sr(N__47303));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__44465),
            .in2(N__44411),
            .in3(N__44438),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__44435),
            .in2(N__44846),
            .in3(N__44414),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__44410),
            .in2(N__44815),
            .in3(N__44384),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__44845),
            .in2(N__44788),
            .in3(N__44819),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__44761),
            .in2(N__44816),
            .in3(N__44792),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__44740),
            .in2(N__44789),
            .in3(N__44765),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__44762),
            .in2(N__44720),
            .in3(N__44744),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__44741),
            .in2(N__44692),
            .in3(N__44723),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47932),
            .ce(N__45377),
            .sr(N__47309));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__44719),
            .in2(N__44659),
            .in3(N__44696),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__44693),
            .in2(N__45139),
            .in3(N__44663),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__45106),
            .in2(N__44660),
            .in3(N__44630),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__45073),
            .in2(N__45140),
            .in3(N__45110),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__45107),
            .in2(N__45038),
            .in3(N__45080),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__45001),
            .in2(N__45077),
            .in3(N__45041),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__45037),
            .in2(N__44971),
            .in3(N__45005),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__45002),
            .in2(N__44932),
            .in3(N__44978),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47924),
            .ce(N__45387),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__44975),
            .in2(N__44878),
            .in3(N__44942),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47917),
            .ce(N__45388),
            .sr(N__47321));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__45436),
            .in2(N__44939),
            .in3(N__44897),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47917),
            .ce(N__45388),
            .sr(N__47321));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__44894),
            .in2(N__44879),
            .in3(N__44849),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47917),
            .ce(N__45388),
            .sr(N__47321));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__45437),
            .in2(N__45419),
            .in3(N__45395),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47917),
            .ce(N__45388),
            .sr(N__47321));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45392),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47917),
            .ce(N__45388),
            .sr(N__47321));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__45338),
            .in2(N__45332),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__45302),
            .in2(_gnd_net_),
            .in3(N__45272),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__45269),
            .in2(N__45263),
            .in3(N__45230),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__45227),
            .in2(_gnd_net_),
            .in3(N__45197),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__45194),
            .in2(_gnd_net_),
            .in3(N__45161),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__45158),
            .in2(_gnd_net_),
            .in3(N__45653),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__45650),
            .in2(_gnd_net_),
            .in3(N__45620),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__45617),
            .in2(_gnd_net_),
            .in3(N__45584),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__45577),
            .in2(_gnd_net_),
            .in3(N__45557),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__45554),
            .in2(_gnd_net_),
            .in3(N__45521),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_20_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__45514),
            .in2(_gnd_net_),
            .in3(N__45494),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_20_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__45487),
            .in2(_gnd_net_),
            .in3(N__45467),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_20_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__45460),
            .in2(_gnd_net_),
            .in3(N__45440),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_20_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__45896),
            .in2(_gnd_net_),
            .in3(N__45866),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_20_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__45859),
            .in2(_gnd_net_),
            .in3(N__45839),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_20_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__45832),
            .in2(_gnd_net_),
            .in3(N__45812),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_21_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__45805),
            .in2(_gnd_net_),
            .in3(N__45785),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_21_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__45778),
            .in2(_gnd_net_),
            .in3(N__45758),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_21_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__45751),
            .in2(_gnd_net_),
            .in3(N__45737),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_18_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_18_21_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_18_21_7  (
            .in0(N__46815),
            .in1(N__46758),
            .in2(_gnd_net_),
            .in3(N__46614),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_18_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_18_22_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_18_22_2  (
            .in0(N__48402),
            .in1(N__48366),
            .in2(N__48055),
            .in3(N__48327),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_20_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_20_15_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_20_15_5  (
            .in0(N__46090),
            .in1(N__46021),
            .in2(N__46468),
            .in3(N__46637),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_2_LC_20_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_2_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_2_LC_20_16_0 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_2_LC_20_16_0  (
            .in0(N__48543),
            .in1(N__46914),
            .in2(N__46734),
            .in3(N__46467),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_18_LC_20_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_18_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_18_LC_20_16_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_18_LC_20_16_1  (
            .in0(N__48154),
            .in1(N__48438),
            .in2(N__46037),
            .in3(N__45983),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_20_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_20_16_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_20_16_2  (
            .in0(N__46030),
            .in1(N__46375),
            .in2(N__45986),
            .in3(N__46647),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_20_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_20_16_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_20_16_3  (
            .in0(_gnd_net_),
            .in1(N__46969),
            .in2(_gnd_net_),
            .in3(N__46591),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_320_4 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_320_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_3_LC_20_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_3_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_3_LC_20_16_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_3_LC_20_16_4  (
            .in0(N__46341),
            .in1(N__46915),
            .in2(N__45977),
            .in3(N__45974),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_20_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_20_16_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_20_16_6  (
            .in0(N__46340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46254),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_20_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_20_16_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_20_16_7  (
            .in0(N__45964),
            .in1(N__48520),
            .in2(N__46699),
            .in3(N__45949),
            .lcout(\delay_measurement_inst.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_20_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_20_17_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_20_17_0  (
            .in0(N__48442),
            .in1(N__46735),
            .in2(N__48147),
            .in3(N__48550),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_20_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_20_17_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_20_17_1  (
            .in0(N__46786),
            .in1(N__45912),
            .in2(N__46850),
            .in3(N__48090),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_331 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_20_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_20_17_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_20_17_2  (
            .in0(N__46272),
            .in1(N__46204),
            .in2(N__46394),
            .in3(N__46391),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_20_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_20_17_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_20_17_3  (
            .in0(N__48252),
            .in1(N__46385),
            .in2(N__46379),
            .in3(N__46363),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_20_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_20_17_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_20_17_4  (
            .in0(N__46273),
            .in1(N__48253),
            .in2(_gnd_net_),
            .in3(N__46206),
            .lcout(\delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_20_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_20_17_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_20_17_6  (
            .in0(N__48091),
            .in1(N__46376),
            .in2(_gnd_net_),
            .in3(N__46205),
            .lcout(\delay_measurement_inst.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_20_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_20_17_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_20_17_7  (
            .in0(N__46274),
            .in1(N__46648),
            .in2(_gnd_net_),
            .in3(N__46364),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_20_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_20_18_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_20_18_0 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_20_18_0  (
            .in0(N__48121),
            .in1(N__46355),
            .in2(N__48257),
            .in3(N__46349),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47933),
            .ce(N__47490),
            .sr(N__47322));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_20_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_20_18_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_20_18_1 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_20_18_1  (
            .in0(N__46275),
            .in1(N__48215),
            .in2(N__46217),
            .in3(N__48122),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47933),
            .ce(N__47490),
            .sr(N__47322));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_20_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_20_18_2 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_20_18_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_20_18_2  (
            .in0(N__46488),
            .in1(N__46536),
            .in2(N__48258),
            .in3(N__46091),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47933),
            .ce(N__47490),
            .sr(N__47322));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_20_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_20_18_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_20_18_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_20_18_3  (
            .in0(N__46534),
            .in1(N__46487),
            .in2(N__46973),
            .in3(N__48216),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47933),
            .ce(N__47490),
            .sr(N__47322));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_20_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_20_18_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_20_18_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_20_18_6  (
            .in0(N__46489),
            .in1(N__46537),
            .in2(N__48259),
            .in3(N__46916),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47933),
            .ce(N__47490),
            .sr(N__47322));
    defparam \delay_measurement_inst.delay_tr_reg_esr_8_LC_20_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_8_LC_20_18_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_8_LC_20_18_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_8_LC_20_18_7  (
            .in0(N__46535),
            .in1(N__48211),
            .in2(_gnd_net_),
            .in3(N__46849),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47933),
            .ce(N__47490),
            .sr(N__47322));
    defparam \delay_measurement_inst.delay_tr_reg_esr_7_LC_20_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_7_LC_20_19_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_7_LC_20_19_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_7_LC_20_19_0  (
            .in0(N__46541),
            .in1(N__48274),
            .in2(_gnd_net_),
            .in3(N__46787),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_20_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_20_19_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_20_19_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_20_19_1  (
            .in0(N__48273),
            .in1(N__46736),
            .in2(_gnd_net_),
            .in3(N__48107),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_20_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_20_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_20_19_3 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_20_19_3  (
            .in0(N__46700),
            .in1(N__48265),
            .in2(_gnd_net_),
            .in3(N__48494),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_20_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_20_19_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_20_19_4 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_20_19_4  (
            .in0(N__46540),
            .in1(N__46499),
            .in2(N__48283),
            .in3(N__46649),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_20_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_20_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_20_19_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_20_19_5  (
            .in0(N__46498),
            .in1(N__46539),
            .in2(N__48284),
            .in3(N__46592),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_20_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_20_19_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_20_19_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_20_19_6  (
            .in0(N__46538),
            .in1(N__46497),
            .in2(N__48282),
            .in3(N__46472),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_20_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_20_19_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_20_19_7 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_20_19_7  (
            .in0(N__48551),
            .in1(N__48266),
            .in2(_gnd_net_),
            .in3(N__48106),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47925),
            .ce(N__47492),
            .sr(N__47327));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_20_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_20_20_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_20_20_0 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_20_20_0  (
            .in0(N__48524),
            .in1(N__48495),
            .in2(_gnd_net_),
            .in3(N__48278),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47918),
            .ce(N__47511),
            .sr(N__47339));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_20_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_20_20_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_20_20_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_20_20_7  (
            .in0(N__48279),
            .in1(N__48443),
            .in2(_gnd_net_),
            .in3(N__48119),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47918),
            .ce(N__47511),
            .sr(N__47339));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_20_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_20_21_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_20_21_2  (
            .in0(N__48388),
            .in1(N__48357),
            .in2(N__48044),
            .in3(N__48318),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_21_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_21_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(N__47459),
            .in2(_gnd_net_),
            .in3(N__48290),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_21_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_21_19_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_21_19_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_21_19_0  (
            .in0(N__48280),
            .in1(N__48155),
            .in2(_gnd_net_),
            .in3(N__48120),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47934),
            .ce(N__47491),
            .sr(N__47340));
endmodule // MAIN
