-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 11 2025 23:51:26

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50432\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50115\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49725\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49601\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10_cascade_\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \N_42_i_i\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_140\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_145\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal un7_start_stop_0_a2 : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_144\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_146\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_71\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_164\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal s4_phy_c : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_204_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_203_i\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal s3_phy_c : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \phase_controller_inst1.N_55_cascade_\ : std_logic;
signal state_ns_i_a2_1 : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \T23_c\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \T45_c\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.N_1326_i\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \phase_controller_inst1.N_55\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.N_54\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \T12_c\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal s1_phy_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_168_i\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_202_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal state_3 : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \T01_c\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_201_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_18_7_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21997\&\N__21990\&\N__21995\&\N__21989\&\N__21996\&\N__21988\&\N__21998\&\N__21985\&\N__21991\&\N__21984\&\N__21992\&\N__21986\&\N__21993\&\N__21987\&\N__21994\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44987\&\N__44984\&'0'&'0'&'0'&\N__44982\&\N__44986\&\N__44983\&\N__44985\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__22010\&\N__22012\&\N__22008\&\N__22011\&\N__22009\&\N__20549\&\N__20565\&\N__20286\&\N__20588\&\N__20273\&\N__20498\&\N__20525\&\N__20443\&\N__20455\&\N__20474\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44879\&\N__44876\&'0'&'0'&'0'&\N__44874\&\N__44878\&\N__44875\&\N__44877\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__28088\,
            RESETB => \N__36362\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__44988\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__44981\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__44925\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__44873\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50430\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50432\,
            DIN => \N__50431\,
            DOUT => \N__50430\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50432\,
            PADOUT => \N__50431\,
            PADIN => \N__50430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50421\,
            DIN => \N__50420\,
            DOUT => \N__50419\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50421\,
            PADOUT => \N__50420\,
            PADIN => \N__50419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__39143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50412\,
            DIN => \N__50411\,
            DOUT => \N__50410\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50412\,
            PADOUT => \N__50411\,
            PADIN => \N__50410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50403\,
            DIN => \N__50402\,
            DOUT => \N__50401\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50403\,
            PADOUT => \N__50402\,
            PADIN => \N__50401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50394\,
            DIN => \N__50393\,
            DOUT => \N__50392\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50394\,
            PADOUT => \N__50393\,
            PADIN => \N__50392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33596\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50385\,
            DIN => \N__50384\,
            DOUT => \N__50383\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50385\,
            PADOUT => \N__50384\,
            PADIN => \N__50383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22196\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50376\,
            DIN => \N__50375\,
            DOUT => \N__50374\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50376\,
            PADOUT => \N__50375\,
            PADIN => \N__50374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50367\,
            DIN => \N__50366\,
            DOUT => \N__50365\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50367\,
            PADOUT => \N__50366\,
            PADIN => \N__50365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35837\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50358\,
            DIN => \N__50357\,
            DOUT => \N__50356\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50358\,
            PADOUT => \N__50357\,
            PADIN => \N__50356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35510\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50349\,
            DIN => \N__50348\,
            DOUT => \N__50347\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50349\,
            PADOUT => \N__50348\,
            PADIN => \N__50347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50340\,
            DIN => \N__50339\,
            DOUT => \N__50338\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50340\,
            PADOUT => \N__50339\,
            PADIN => \N__50338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50331\,
            DIN => \N__50330\,
            DOUT => \N__50329\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50331\,
            PADOUT => \N__50330\,
            PADIN => \N__50329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25445\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50322\,
            DIN => \N__50321\,
            DOUT => \N__50320\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50322\,
            PADOUT => \N__50321\,
            PADIN => \N__50320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50313\,
            DIN => \N__50312\,
            DOUT => \N__50311\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50313\,
            PADOUT => \N__50312\,
            PADIN => \N__50311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28109\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50304\,
            DIN => \N__50303\,
            DOUT => \N__50302\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50304\,
            PADOUT => \N__50303\,
            PADIN => \N__50302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33551\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50295\,
            DIN => \N__50294\,
            DOUT => \N__50293\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50295\,
            PADOUT => \N__50294\,
            PADIN => \N__50293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50286\,
            DIN => \N__50285\,
            DOUT => \N__50284\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50286\,
            PADOUT => \N__50285\,
            PADIN => \N__50284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11929\ : InMux
    port map (
            O => \N__50267\,
            I => \N__50264\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__50264\,
            I => \N__50261\
        );

    \I__11927\ : Span4Mux_v
    port map (
            O => \N__50261\,
            I => \N__50255\
        );

    \I__11926\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50252\
        );

    \I__11925\ : InMux
    port map (
            O => \N__50259\,
            I => \N__50249\
        );

    \I__11924\ : InMux
    port map (
            O => \N__50258\,
            I => \N__50246\
        );

    \I__11923\ : Odrv4
    port map (
            O => \N__50255\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__50252\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__50249\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11920\ : LocalMux
    port map (
            O => \N__50246\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__11919\ : InMux
    port map (
            O => \N__50237\,
            I => \N__50232\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50236\,
            I => \N__50229\
        );

    \I__11917\ : InMux
    port map (
            O => \N__50235\,
            I => \N__50226\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__50232\,
            I => \N__50223\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__50229\,
            I => \N__50220\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__50226\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11913\ : Odrv4
    port map (
            O => \N__50223\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11912\ : Odrv4
    port map (
            O => \N__50220\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__11911\ : CascadeMux
    port map (
            O => \N__50213\,
            I => \N__50209\
        );

    \I__11910\ : CascadeMux
    port map (
            O => \N__50212\,
            I => \N__50206\
        );

    \I__11909\ : InMux
    port map (
            O => \N__50209\,
            I => \N__50201\
        );

    \I__11908\ : InMux
    port map (
            O => \N__50206\,
            I => \N__50201\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__50201\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__11906\ : InMux
    port map (
            O => \N__50198\,
            I => \N__50194\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50197\,
            I => \N__50190\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__50194\,
            I => \N__50187\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50193\,
            I => \N__50184\
        );

    \I__11902\ : LocalMux
    port map (
            O => \N__50190\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11901\ : Odrv12
    port map (
            O => \N__50187\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__50184\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11899\ : InMux
    port map (
            O => \N__50177\,
            I => \N__50174\
        );

    \I__11898\ : LocalMux
    port map (
            O => \N__50174\,
            I => \N__50169\
        );

    \I__11897\ : InMux
    port map (
            O => \N__50173\,
            I => \N__50166\
        );

    \I__11896\ : InMux
    port map (
            O => \N__50172\,
            I => \N__50163\
        );

    \I__11895\ : Span4Mux_v
    port map (
            O => \N__50169\,
            I => \N__50157\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__50166\,
            I => \N__50157\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__50163\,
            I => \N__50154\
        );

    \I__11892\ : InMux
    port map (
            O => \N__50162\,
            I => \N__50151\
        );

    \I__11891\ : Odrv4
    port map (
            O => \N__50157\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__11890\ : Odrv4
    port map (
            O => \N__50154\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__50151\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__11888\ : InMux
    port map (
            O => \N__50144\,
            I => \N__50138\
        );

    \I__11887\ : InMux
    port map (
            O => \N__50143\,
            I => \N__50138\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__50138\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__11885\ : InMux
    port map (
            O => \N__50135\,
            I => \N__50129\
        );

    \I__11884\ : InMux
    port map (
            O => \N__50134\,
            I => \N__50126\
        );

    \I__11883\ : InMux
    port map (
            O => \N__50133\,
            I => \N__50121\
        );

    \I__11882\ : InMux
    port map (
            O => \N__50132\,
            I => \N__50121\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__50129\,
            I => \N__50118\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__50126\,
            I => \N__50115\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__50121\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__11878\ : Odrv12
    port map (
            O => \N__50118\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__11877\ : Odrv4
    port map (
            O => \N__50115\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__11876\ : CascadeMux
    port map (
            O => \N__50108\,
            I => \N__50105\
        );

    \I__11875\ : InMux
    port map (
            O => \N__50105\,
            I => \N__50102\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__50102\,
            I => \N__50095\
        );

    \I__11873\ : InMux
    port map (
            O => \N__50101\,
            I => \N__50092\
        );

    \I__11872\ : InMux
    port map (
            O => \N__50100\,
            I => \N__50089\
        );

    \I__11871\ : InMux
    port map (
            O => \N__50099\,
            I => \N__50084\
        );

    \I__11870\ : InMux
    port map (
            O => \N__50098\,
            I => \N__50084\
        );

    \I__11869\ : Span4Mux_v
    port map (
            O => \N__50095\,
            I => \N__50079\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__50092\,
            I => \N__50079\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__50089\,
            I => \N__50074\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__50084\,
            I => \N__50074\
        );

    \I__11865\ : Span4Mux_h
    port map (
            O => \N__50079\,
            I => \N__50071\
        );

    \I__11864\ : Odrv12
    port map (
            O => \N__50074\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__11863\ : Odrv4
    port map (
            O => \N__50071\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__11862\ : CEMux
    port map (
            O => \N__50066\,
            I => \N__50063\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__50063\,
            I => \N__50059\
        );

    \I__11860\ : CEMux
    port map (
            O => \N__50062\,
            I => \N__50056\
        );

    \I__11859\ : Span4Mux_v
    port map (
            O => \N__50059\,
            I => \N__50042\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__50056\,
            I => \N__50042\
        );

    \I__11857\ : InMux
    port map (
            O => \N__50055\,
            I => \N__50035\
        );

    \I__11856\ : InMux
    port map (
            O => \N__50054\,
            I => \N__50035\
        );

    \I__11855\ : InMux
    port map (
            O => \N__50053\,
            I => \N__50035\
        );

    \I__11854\ : InMux
    port map (
            O => \N__50052\,
            I => \N__50028\
        );

    \I__11853\ : InMux
    port map (
            O => \N__50051\,
            I => \N__50018\
        );

    \I__11852\ : InMux
    port map (
            O => \N__50050\,
            I => \N__50018\
        );

    \I__11851\ : InMux
    port map (
            O => \N__50049\,
            I => \N__50018\
        );

    \I__11850\ : InMux
    port map (
            O => \N__50048\,
            I => \N__50018\
        );

    \I__11849\ : CEMux
    port map (
            O => \N__50047\,
            I => \N__50015\
        );

    \I__11848\ : Span4Mux_h
    port map (
            O => \N__50042\,
            I => \N__50010\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__50035\,
            I => \N__50010\
        );

    \I__11846\ : CEMux
    port map (
            O => \N__50034\,
            I => \N__50007\
        );

    \I__11845\ : CEMux
    port map (
            O => \N__50033\,
            I => \N__50002\
        );

    \I__11844\ : CEMux
    port map (
            O => \N__50032\,
            I => \N__49995\
        );

    \I__11843\ : CEMux
    port map (
            O => \N__50031\,
            I => \N__49991\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__50028\,
            I => \N__49987\
        );

    \I__11841\ : CEMux
    port map (
            O => \N__50027\,
            I => \N__49984\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__50018\,
            I => \N__49970\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__50015\,
            I => \N__49970\
        );

    \I__11838\ : Span4Mux_v
    port map (
            O => \N__50010\,
            I => \N__49965\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__50007\,
            I => \N__49965\
        );

    \I__11836\ : CEMux
    port map (
            O => \N__50006\,
            I => \N__49949\
        );

    \I__11835\ : CEMux
    port map (
            O => \N__50005\,
            I => \N__49946\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__50002\,
            I => \N__49943\
        );

    \I__11833\ : InMux
    port map (
            O => \N__50001\,
            I => \N__49934\
        );

    \I__11832\ : InMux
    port map (
            O => \N__50000\,
            I => \N__49934\
        );

    \I__11831\ : InMux
    port map (
            O => \N__49999\,
            I => \N__49934\
        );

    \I__11830\ : InMux
    port map (
            O => \N__49998\,
            I => \N__49934\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__49995\,
            I => \N__49931\
        );

    \I__11828\ : CEMux
    port map (
            O => \N__49994\,
            I => \N__49928\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__49991\,
            I => \N__49925\
        );

    \I__11826\ : CEMux
    port map (
            O => \N__49990\,
            I => \N__49922\
        );

    \I__11825\ : Span4Mux_v
    port map (
            O => \N__49987\,
            I => \N__49917\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__49984\,
            I => \N__49917\
        );

    \I__11823\ : CEMux
    port map (
            O => \N__49983\,
            I => \N__49914\
        );

    \I__11822\ : CEMux
    port map (
            O => \N__49982\,
            I => \N__49911\
        );

    \I__11821\ : InMux
    port map (
            O => \N__49981\,
            I => \N__49902\
        );

    \I__11820\ : InMux
    port map (
            O => \N__49980\,
            I => \N__49902\
        );

    \I__11819\ : InMux
    port map (
            O => \N__49979\,
            I => \N__49902\
        );

    \I__11818\ : InMux
    port map (
            O => \N__49978\,
            I => \N__49902\
        );

    \I__11817\ : InMux
    port map (
            O => \N__49977\,
            I => \N__49895\
        );

    \I__11816\ : InMux
    port map (
            O => \N__49976\,
            I => \N__49895\
        );

    \I__11815\ : InMux
    port map (
            O => \N__49975\,
            I => \N__49895\
        );

    \I__11814\ : Span4Mux_v
    port map (
            O => \N__49970\,
            I => \N__49890\
        );

    \I__11813\ : Span4Mux_v
    port map (
            O => \N__49965\,
            I => \N__49890\
        );

    \I__11812\ : InMux
    port map (
            O => \N__49964\,
            I => \N__49881\
        );

    \I__11811\ : InMux
    port map (
            O => \N__49963\,
            I => \N__49881\
        );

    \I__11810\ : InMux
    port map (
            O => \N__49962\,
            I => \N__49881\
        );

    \I__11809\ : InMux
    port map (
            O => \N__49961\,
            I => \N__49881\
        );

    \I__11808\ : InMux
    port map (
            O => \N__49960\,
            I => \N__49872\
        );

    \I__11807\ : InMux
    port map (
            O => \N__49959\,
            I => \N__49872\
        );

    \I__11806\ : InMux
    port map (
            O => \N__49958\,
            I => \N__49872\
        );

    \I__11805\ : InMux
    port map (
            O => \N__49957\,
            I => \N__49872\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49956\,
            I => \N__49863\
        );

    \I__11803\ : InMux
    port map (
            O => \N__49955\,
            I => \N__49863\
        );

    \I__11802\ : InMux
    port map (
            O => \N__49954\,
            I => \N__49863\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49953\,
            I => \N__49863\
        );

    \I__11800\ : CEMux
    port map (
            O => \N__49952\,
            I => \N__49860\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__49949\,
            I => \N__49855\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__49946\,
            I => \N__49855\
        );

    \I__11797\ : Span4Mux_h
    port map (
            O => \N__49943\,
            I => \N__49852\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__49934\,
            I => \N__49849\
        );

    \I__11795\ : Span4Mux_h
    port map (
            O => \N__49931\,
            I => \N__49846\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__49928\,
            I => \N__49837\
        );

    \I__11793\ : Span4Mux_h
    port map (
            O => \N__49925\,
            I => \N__49837\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__49922\,
            I => \N__49837\
        );

    \I__11791\ : Span4Mux_h
    port map (
            O => \N__49917\,
            I => \N__49837\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__49914\,
            I => \N__49834\
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__49911\,
            I => \N__49831\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__49902\,
            I => \N__49818\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__49895\,
            I => \N__49818\
        );

    \I__11786\ : Span4Mux_h
    port map (
            O => \N__49890\,
            I => \N__49818\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__49881\,
            I => \N__49818\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__49872\,
            I => \N__49818\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__49863\,
            I => \N__49818\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49860\,
            I => \N__49815\
        );

    \I__11781\ : Span4Mux_h
    port map (
            O => \N__49855\,
            I => \N__49810\
        );

    \I__11780\ : Span4Mux_h
    port map (
            O => \N__49852\,
            I => \N__49810\
        );

    \I__11779\ : Span4Mux_h
    port map (
            O => \N__49849\,
            I => \N__49801\
        );

    \I__11778\ : Span4Mux_h
    port map (
            O => \N__49846\,
            I => \N__49801\
        );

    \I__11777\ : Span4Mux_h
    port map (
            O => \N__49837\,
            I => \N__49801\
        );

    \I__11776\ : Span4Mux_h
    port map (
            O => \N__49834\,
            I => \N__49801\
        );

    \I__11775\ : Span12Mux_h
    port map (
            O => \N__49831\,
            I => \N__49798\
        );

    \I__11774\ : Span4Mux_v
    port map (
            O => \N__49818\,
            I => \N__49795\
        );

    \I__11773\ : Span4Mux_h
    port map (
            O => \N__49815\,
            I => \N__49790\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__49810\,
            I => \N__49790\
        );

    \I__11771\ : Span4Mux_v
    port map (
            O => \N__49801\,
            I => \N__49787\
        );

    \I__11770\ : Odrv12
    port map (
            O => \N__49798\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11769\ : Odrv4
    port map (
            O => \N__49795\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11768\ : Odrv4
    port map (
            O => \N__49790\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11767\ : Odrv4
    port map (
            O => \N__49787\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11766\ : InMux
    port map (
            O => \N__49778\,
            I => \N__49774\
        );

    \I__11765\ : CascadeMux
    port map (
            O => \N__49777\,
            I => \N__49770\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__49774\,
            I => \N__49766\
        );

    \I__11763\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49763\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49770\,
            I => \N__49760\
        );

    \I__11761\ : InMux
    port map (
            O => \N__49769\,
            I => \N__49757\
        );

    \I__11760\ : Span4Mux_h
    port map (
            O => \N__49766\,
            I => \N__49754\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__49763\,
            I => \N__49749\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__49760\,
            I => \N__49749\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__49757\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__11756\ : Odrv4
    port map (
            O => \N__49754\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__11755\ : Odrv12
    port map (
            O => \N__49749\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49738\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49741\,
            I => \N__49735\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__49738\,
            I => \N__49731\
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__49735\,
            I => \N__49728\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49734\,
            I => \N__49725\
        );

    \I__11749\ : Span4Mux_h
    port map (
            O => \N__49731\,
            I => \N__49720\
        );

    \I__11748\ : Span4Mux_v
    port map (
            O => \N__49728\,
            I => \N__49720\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__49725\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__11746\ : Odrv4
    port map (
            O => \N__49720\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__11745\ : InMux
    port map (
            O => \N__49715\,
            I => \N__49710\
        );

    \I__11744\ : InMux
    port map (
            O => \N__49714\,
            I => \N__49706\
        );

    \I__11743\ : InMux
    port map (
            O => \N__49713\,
            I => \N__49703\
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__49710\,
            I => \N__49700\
        );

    \I__11741\ : InMux
    port map (
            O => \N__49709\,
            I => \N__49697\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__49706\,
            I => \N__49694\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__49703\,
            I => \N__49691\
        );

    \I__11738\ : Span4Mux_v
    port map (
            O => \N__49700\,
            I => \N__49688\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__49697\,
            I => \N__49685\
        );

    \I__11736\ : Span4Mux_v
    port map (
            O => \N__49694\,
            I => \N__49682\
        );

    \I__11735\ : Span12Mux_s9_h
    port map (
            O => \N__49691\,
            I => \N__49679\
        );

    \I__11734\ : Span4Mux_h
    port map (
            O => \N__49688\,
            I => \N__49674\
        );

    \I__11733\ : Span4Mux_h
    port map (
            O => \N__49685\,
            I => \N__49674\
        );

    \I__11732\ : Odrv4
    port map (
            O => \N__49682\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11731\ : Odrv12
    port map (
            O => \N__49679\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11730\ : Odrv4
    port map (
            O => \N__49674\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49667\,
            I => \N__49663\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49666\,
            I => \N__49660\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__49663\,
            I => \N__49656\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__49660\,
            I => \N__49653\
        );

    \I__11725\ : InMux
    port map (
            O => \N__49659\,
            I => \N__49650\
        );

    \I__11724\ : Span4Mux_v
    port map (
            O => \N__49656\,
            I => \N__49645\
        );

    \I__11723\ : Span4Mux_h
    port map (
            O => \N__49653\,
            I => \N__49645\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__49650\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__11721\ : Odrv4
    port map (
            O => \N__49645\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__11720\ : InMux
    port map (
            O => \N__49640\,
            I => \N__49632\
        );

    \I__11719\ : InMux
    port map (
            O => \N__49639\,
            I => \N__49620\
        );

    \I__11718\ : InMux
    port map (
            O => \N__49638\,
            I => \N__49604\
        );

    \I__11717\ : InMux
    port map (
            O => \N__49637\,
            I => \N__49604\
        );

    \I__11716\ : InMux
    port map (
            O => \N__49636\,
            I => \N__49604\
        );

    \I__11715\ : InMux
    port map (
            O => \N__49635\,
            I => \N__49604\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__49632\,
            I => \N__49601\
        );

    \I__11713\ : InMux
    port map (
            O => \N__49631\,
            I => \N__49594\
        );

    \I__11712\ : InMux
    port map (
            O => \N__49630\,
            I => \N__49594\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49629\,
            I => \N__49594\
        );

    \I__11710\ : InMux
    port map (
            O => \N__49628\,
            I => \N__49556\
        );

    \I__11709\ : InMux
    port map (
            O => \N__49627\,
            I => \N__49556\
        );

    \I__11708\ : InMux
    port map (
            O => \N__49626\,
            I => \N__49556\
        );

    \I__11707\ : InMux
    port map (
            O => \N__49625\,
            I => \N__49556\
        );

    \I__11706\ : InMux
    port map (
            O => \N__49624\,
            I => \N__49556\
        );

    \I__11705\ : CascadeMux
    port map (
            O => \N__49623\,
            I => \N__49551\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__49620\,
            I => \N__49543\
        );

    \I__11703\ : InMux
    port map (
            O => \N__49619\,
            I => \N__49538\
        );

    \I__11702\ : InMux
    port map (
            O => \N__49618\,
            I => \N__49538\
        );

    \I__11701\ : InMux
    port map (
            O => \N__49617\,
            I => \N__49535\
        );

    \I__11700\ : InMux
    port map (
            O => \N__49616\,
            I => \N__49527\
        );

    \I__11699\ : InMux
    port map (
            O => \N__49615\,
            I => \N__49520\
        );

    \I__11698\ : InMux
    port map (
            O => \N__49614\,
            I => \N__49520\
        );

    \I__11697\ : InMux
    port map (
            O => \N__49613\,
            I => \N__49520\
        );

    \I__11696\ : LocalMux
    port map (
            O => \N__49604\,
            I => \N__49517\
        );

    \I__11695\ : Span4Mux_h
    port map (
            O => \N__49601\,
            I => \N__49512\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__49594\,
            I => \N__49512\
        );

    \I__11693\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49509\
        );

    \I__11692\ : InMux
    port map (
            O => \N__49592\,
            I => \N__49498\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49591\,
            I => \N__49498\
        );

    \I__11690\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49498\
        );

    \I__11689\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49498\
        );

    \I__11688\ : InMux
    port map (
            O => \N__49588\,
            I => \N__49498\
        );

    \I__11687\ : InMux
    port map (
            O => \N__49587\,
            I => \N__49489\
        );

    \I__11686\ : InMux
    port map (
            O => \N__49586\,
            I => \N__49489\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49585\,
            I => \N__49489\
        );

    \I__11684\ : InMux
    port map (
            O => \N__49584\,
            I => \N__49489\
        );

    \I__11683\ : InMux
    port map (
            O => \N__49583\,
            I => \N__49482\
        );

    \I__11682\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49482\
        );

    \I__11681\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49482\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49476\
        );

    \I__11679\ : CascadeMux
    port map (
            O => \N__49579\,
            I => \N__49473\
        );

    \I__11678\ : CascadeMux
    port map (
            O => \N__49578\,
            I => \N__49470\
        );

    \I__11677\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49466\
        );

    \I__11676\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49459\
        );

    \I__11675\ : InMux
    port map (
            O => \N__49575\,
            I => \N__49459\
        );

    \I__11674\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49459\
        );

    \I__11673\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49447\
        );

    \I__11672\ : InMux
    port map (
            O => \N__49572\,
            I => \N__49447\
        );

    \I__11671\ : InMux
    port map (
            O => \N__49571\,
            I => \N__49436\
        );

    \I__11670\ : InMux
    port map (
            O => \N__49570\,
            I => \N__49436\
        );

    \I__11669\ : InMux
    port map (
            O => \N__49569\,
            I => \N__49436\
        );

    \I__11668\ : InMux
    port map (
            O => \N__49568\,
            I => \N__49436\
        );

    \I__11667\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49436\
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__49556\,
            I => \N__49433\
        );

    \I__11665\ : InMux
    port map (
            O => \N__49555\,
            I => \N__49430\
        );

    \I__11664\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49426\
        );

    \I__11663\ : InMux
    port map (
            O => \N__49551\,
            I => \N__49415\
        );

    \I__11662\ : InMux
    port map (
            O => \N__49550\,
            I => \N__49408\
        );

    \I__11661\ : InMux
    port map (
            O => \N__49549\,
            I => \N__49408\
        );

    \I__11660\ : InMux
    port map (
            O => \N__49548\,
            I => \N__49408\
        );

    \I__11659\ : InMux
    port map (
            O => \N__49547\,
            I => \N__49403\
        );

    \I__11658\ : InMux
    port map (
            O => \N__49546\,
            I => \N__49403\
        );

    \I__11657\ : Span4Mux_v
    port map (
            O => \N__49543\,
            I => \N__49400\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__49538\,
            I => \N__49395\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__49535\,
            I => \N__49395\
        );

    \I__11654\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49392\
        );

    \I__11653\ : InMux
    port map (
            O => \N__49533\,
            I => \N__49383\
        );

    \I__11652\ : InMux
    port map (
            O => \N__49532\,
            I => \N__49383\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49531\,
            I => \N__49383\
        );

    \I__11650\ : InMux
    port map (
            O => \N__49530\,
            I => \N__49383\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__49527\,
            I => \N__49372\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__49520\,
            I => \N__49372\
        );

    \I__11647\ : Span4Mux_v
    port map (
            O => \N__49517\,
            I => \N__49372\
        );

    \I__11646\ : Span4Mux_v
    port map (
            O => \N__49512\,
            I => \N__49372\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__49509\,
            I => \N__49372\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__49498\,
            I => \N__49367\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__49489\,
            I => \N__49367\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__49482\,
            I => \N__49364\
        );

    \I__11641\ : InMux
    port map (
            O => \N__49481\,
            I => \N__49357\
        );

    \I__11640\ : InMux
    port map (
            O => \N__49480\,
            I => \N__49357\
        );

    \I__11639\ : InMux
    port map (
            O => \N__49479\,
            I => \N__49357\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__49476\,
            I => \N__49354\
        );

    \I__11637\ : InMux
    port map (
            O => \N__49473\,
            I => \N__49343\
        );

    \I__11636\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49343\
        );

    \I__11635\ : InMux
    port map (
            O => \N__49469\,
            I => \N__49343\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__49466\,
            I => \N__49340\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__49459\,
            I => \N__49337\
        );

    \I__11632\ : InMux
    port map (
            O => \N__49458\,
            I => \N__49329\
        );

    \I__11631\ : InMux
    port map (
            O => \N__49457\,
            I => \N__49329\
        );

    \I__11630\ : InMux
    port map (
            O => \N__49456\,
            I => \N__49322\
        );

    \I__11629\ : InMux
    port map (
            O => \N__49455\,
            I => \N__49322\
        );

    \I__11628\ : InMux
    port map (
            O => \N__49454\,
            I => \N__49322\
        );

    \I__11627\ : InMux
    port map (
            O => \N__49453\,
            I => \N__49313\
        );

    \I__11626\ : InMux
    port map (
            O => \N__49452\,
            I => \N__49313\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__49447\,
            I => \N__49304\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__49436\,
            I => \N__49304\
        );

    \I__11623\ : Sp12to4
    port map (
            O => \N__49433\,
            I => \N__49304\
        );

    \I__11622\ : LocalMux
    port map (
            O => \N__49430\,
            I => \N__49304\
        );

    \I__11621\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49301\
        );

    \I__11620\ : LocalMux
    port map (
            O => \N__49426\,
            I => \N__49298\
        );

    \I__11619\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49295\
        );

    \I__11618\ : InMux
    port map (
            O => \N__49424\,
            I => \N__49288\
        );

    \I__11617\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49288\
        );

    \I__11616\ : InMux
    port map (
            O => \N__49422\,
            I => \N__49288\
        );

    \I__11615\ : InMux
    port map (
            O => \N__49421\,
            I => \N__49281\
        );

    \I__11614\ : InMux
    port map (
            O => \N__49420\,
            I => \N__49281\
        );

    \I__11613\ : InMux
    port map (
            O => \N__49419\,
            I => \N__49281\
        );

    \I__11612\ : InMux
    port map (
            O => \N__49418\,
            I => \N__49278\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__49415\,
            I => \N__49267\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__49408\,
            I => \N__49267\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__49403\,
            I => \N__49267\
        );

    \I__11608\ : Span4Mux_h
    port map (
            O => \N__49400\,
            I => \N__49267\
        );

    \I__11607\ : Span4Mux_h
    port map (
            O => \N__49395\,
            I => \N__49267\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__49392\,
            I => \N__49264\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__49383\,
            I => \N__49257\
        );

    \I__11604\ : Span4Mux_v
    port map (
            O => \N__49372\,
            I => \N__49257\
        );

    \I__11603\ : Span4Mux_v
    port map (
            O => \N__49367\,
            I => \N__49257\
        );

    \I__11602\ : Span4Mux_h
    port map (
            O => \N__49364\,
            I => \N__49250\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__49357\,
            I => \N__49250\
        );

    \I__11600\ : Span4Mux_v
    port map (
            O => \N__49354\,
            I => \N__49250\
        );

    \I__11599\ : InMux
    port map (
            O => \N__49353\,
            I => \N__49247\
        );

    \I__11598\ : InMux
    port map (
            O => \N__49352\,
            I => \N__49242\
        );

    \I__11597\ : InMux
    port map (
            O => \N__49351\,
            I => \N__49242\
        );

    \I__11596\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49239\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__49343\,
            I => \N__49232\
        );

    \I__11594\ : Span4Mux_h
    port map (
            O => \N__49340\,
            I => \N__49232\
        );

    \I__11593\ : Span4Mux_h
    port map (
            O => \N__49337\,
            I => \N__49232\
        );

    \I__11592\ : InMux
    port map (
            O => \N__49336\,
            I => \N__49229\
        );

    \I__11591\ : InMux
    port map (
            O => \N__49335\,
            I => \N__49224\
        );

    \I__11590\ : InMux
    port map (
            O => \N__49334\,
            I => \N__49224\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__49329\,
            I => \N__49219\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__49322\,
            I => \N__49219\
        );

    \I__11587\ : InMux
    port map (
            O => \N__49321\,
            I => \N__49210\
        );

    \I__11586\ : InMux
    port map (
            O => \N__49320\,
            I => \N__49210\
        );

    \I__11585\ : InMux
    port map (
            O => \N__49319\,
            I => \N__49210\
        );

    \I__11584\ : InMux
    port map (
            O => \N__49318\,
            I => \N__49210\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__49313\,
            I => \N__49203\
        );

    \I__11582\ : Span12Mux_h
    port map (
            O => \N__49304\,
            I => \N__49203\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__49301\,
            I => \N__49203\
        );

    \I__11580\ : Span4Mux_v
    port map (
            O => \N__49298\,
            I => \N__49196\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__49295\,
            I => \N__49196\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__49288\,
            I => \N__49196\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__49281\,
            I => \N__49189\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__49278\,
            I => \N__49189\
        );

    \I__11575\ : Span4Mux_h
    port map (
            O => \N__49267\,
            I => \N__49189\
        );

    \I__11574\ : Span4Mux_h
    port map (
            O => \N__49264\,
            I => \N__49182\
        );

    \I__11573\ : Span4Mux_h
    port map (
            O => \N__49257\,
            I => \N__49182\
        );

    \I__11572\ : Span4Mux_v
    port map (
            O => \N__49250\,
            I => \N__49182\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__49247\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__49242\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__49239\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11568\ : Odrv4
    port map (
            O => \N__49232\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__49229\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__49224\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11565\ : Odrv12
    port map (
            O => \N__49219\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__49210\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11563\ : Odrv12
    port map (
            O => \N__49203\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11562\ : Odrv4
    port map (
            O => \N__49196\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11561\ : Odrv4
    port map (
            O => \N__49189\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11560\ : Odrv4
    port map (
            O => \N__49182\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49157\,
            I => \N__49154\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__49154\,
            I => \N__49151\
        );

    \I__11557\ : Odrv12
    port map (
            O => \N__49151\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__11556\ : ClkMux
    port map (
            O => \N__49148\,
            I => \N__48725\
        );

    \I__11555\ : ClkMux
    port map (
            O => \N__49147\,
            I => \N__48725\
        );

    \I__11554\ : ClkMux
    port map (
            O => \N__49146\,
            I => \N__48725\
        );

    \I__11553\ : ClkMux
    port map (
            O => \N__49145\,
            I => \N__48725\
        );

    \I__11552\ : ClkMux
    port map (
            O => \N__49144\,
            I => \N__48725\
        );

    \I__11551\ : ClkMux
    port map (
            O => \N__49143\,
            I => \N__48725\
        );

    \I__11550\ : ClkMux
    port map (
            O => \N__49142\,
            I => \N__48725\
        );

    \I__11549\ : ClkMux
    port map (
            O => \N__49141\,
            I => \N__48725\
        );

    \I__11548\ : ClkMux
    port map (
            O => \N__49140\,
            I => \N__48725\
        );

    \I__11547\ : ClkMux
    port map (
            O => \N__49139\,
            I => \N__48725\
        );

    \I__11546\ : ClkMux
    port map (
            O => \N__49138\,
            I => \N__48725\
        );

    \I__11545\ : ClkMux
    port map (
            O => \N__49137\,
            I => \N__48725\
        );

    \I__11544\ : ClkMux
    port map (
            O => \N__49136\,
            I => \N__48725\
        );

    \I__11543\ : ClkMux
    port map (
            O => \N__49135\,
            I => \N__48725\
        );

    \I__11542\ : ClkMux
    port map (
            O => \N__49134\,
            I => \N__48725\
        );

    \I__11541\ : ClkMux
    port map (
            O => \N__49133\,
            I => \N__48725\
        );

    \I__11540\ : ClkMux
    port map (
            O => \N__49132\,
            I => \N__48725\
        );

    \I__11539\ : ClkMux
    port map (
            O => \N__49131\,
            I => \N__48725\
        );

    \I__11538\ : ClkMux
    port map (
            O => \N__49130\,
            I => \N__48725\
        );

    \I__11537\ : ClkMux
    port map (
            O => \N__49129\,
            I => \N__48725\
        );

    \I__11536\ : ClkMux
    port map (
            O => \N__49128\,
            I => \N__48725\
        );

    \I__11535\ : ClkMux
    port map (
            O => \N__49127\,
            I => \N__48725\
        );

    \I__11534\ : ClkMux
    port map (
            O => \N__49126\,
            I => \N__48725\
        );

    \I__11533\ : ClkMux
    port map (
            O => \N__49125\,
            I => \N__48725\
        );

    \I__11532\ : ClkMux
    port map (
            O => \N__49124\,
            I => \N__48725\
        );

    \I__11531\ : ClkMux
    port map (
            O => \N__49123\,
            I => \N__48725\
        );

    \I__11530\ : ClkMux
    port map (
            O => \N__49122\,
            I => \N__48725\
        );

    \I__11529\ : ClkMux
    port map (
            O => \N__49121\,
            I => \N__48725\
        );

    \I__11528\ : ClkMux
    port map (
            O => \N__49120\,
            I => \N__48725\
        );

    \I__11527\ : ClkMux
    port map (
            O => \N__49119\,
            I => \N__48725\
        );

    \I__11526\ : ClkMux
    port map (
            O => \N__49118\,
            I => \N__48725\
        );

    \I__11525\ : ClkMux
    port map (
            O => \N__49117\,
            I => \N__48725\
        );

    \I__11524\ : ClkMux
    port map (
            O => \N__49116\,
            I => \N__48725\
        );

    \I__11523\ : ClkMux
    port map (
            O => \N__49115\,
            I => \N__48725\
        );

    \I__11522\ : ClkMux
    port map (
            O => \N__49114\,
            I => \N__48725\
        );

    \I__11521\ : ClkMux
    port map (
            O => \N__49113\,
            I => \N__48725\
        );

    \I__11520\ : ClkMux
    port map (
            O => \N__49112\,
            I => \N__48725\
        );

    \I__11519\ : ClkMux
    port map (
            O => \N__49111\,
            I => \N__48725\
        );

    \I__11518\ : ClkMux
    port map (
            O => \N__49110\,
            I => \N__48725\
        );

    \I__11517\ : ClkMux
    port map (
            O => \N__49109\,
            I => \N__48725\
        );

    \I__11516\ : ClkMux
    port map (
            O => \N__49108\,
            I => \N__48725\
        );

    \I__11515\ : ClkMux
    port map (
            O => \N__49107\,
            I => \N__48725\
        );

    \I__11514\ : ClkMux
    port map (
            O => \N__49106\,
            I => \N__48725\
        );

    \I__11513\ : ClkMux
    port map (
            O => \N__49105\,
            I => \N__48725\
        );

    \I__11512\ : ClkMux
    port map (
            O => \N__49104\,
            I => \N__48725\
        );

    \I__11511\ : ClkMux
    port map (
            O => \N__49103\,
            I => \N__48725\
        );

    \I__11510\ : ClkMux
    port map (
            O => \N__49102\,
            I => \N__48725\
        );

    \I__11509\ : ClkMux
    port map (
            O => \N__49101\,
            I => \N__48725\
        );

    \I__11508\ : ClkMux
    port map (
            O => \N__49100\,
            I => \N__48725\
        );

    \I__11507\ : ClkMux
    port map (
            O => \N__49099\,
            I => \N__48725\
        );

    \I__11506\ : ClkMux
    port map (
            O => \N__49098\,
            I => \N__48725\
        );

    \I__11505\ : ClkMux
    port map (
            O => \N__49097\,
            I => \N__48725\
        );

    \I__11504\ : ClkMux
    port map (
            O => \N__49096\,
            I => \N__48725\
        );

    \I__11503\ : ClkMux
    port map (
            O => \N__49095\,
            I => \N__48725\
        );

    \I__11502\ : ClkMux
    port map (
            O => \N__49094\,
            I => \N__48725\
        );

    \I__11501\ : ClkMux
    port map (
            O => \N__49093\,
            I => \N__48725\
        );

    \I__11500\ : ClkMux
    port map (
            O => \N__49092\,
            I => \N__48725\
        );

    \I__11499\ : ClkMux
    port map (
            O => \N__49091\,
            I => \N__48725\
        );

    \I__11498\ : ClkMux
    port map (
            O => \N__49090\,
            I => \N__48725\
        );

    \I__11497\ : ClkMux
    port map (
            O => \N__49089\,
            I => \N__48725\
        );

    \I__11496\ : ClkMux
    port map (
            O => \N__49088\,
            I => \N__48725\
        );

    \I__11495\ : ClkMux
    port map (
            O => \N__49087\,
            I => \N__48725\
        );

    \I__11494\ : ClkMux
    port map (
            O => \N__49086\,
            I => \N__48725\
        );

    \I__11493\ : ClkMux
    port map (
            O => \N__49085\,
            I => \N__48725\
        );

    \I__11492\ : ClkMux
    port map (
            O => \N__49084\,
            I => \N__48725\
        );

    \I__11491\ : ClkMux
    port map (
            O => \N__49083\,
            I => \N__48725\
        );

    \I__11490\ : ClkMux
    port map (
            O => \N__49082\,
            I => \N__48725\
        );

    \I__11489\ : ClkMux
    port map (
            O => \N__49081\,
            I => \N__48725\
        );

    \I__11488\ : ClkMux
    port map (
            O => \N__49080\,
            I => \N__48725\
        );

    \I__11487\ : ClkMux
    port map (
            O => \N__49079\,
            I => \N__48725\
        );

    \I__11486\ : ClkMux
    port map (
            O => \N__49078\,
            I => \N__48725\
        );

    \I__11485\ : ClkMux
    port map (
            O => \N__49077\,
            I => \N__48725\
        );

    \I__11484\ : ClkMux
    port map (
            O => \N__49076\,
            I => \N__48725\
        );

    \I__11483\ : ClkMux
    port map (
            O => \N__49075\,
            I => \N__48725\
        );

    \I__11482\ : ClkMux
    port map (
            O => \N__49074\,
            I => \N__48725\
        );

    \I__11481\ : ClkMux
    port map (
            O => \N__49073\,
            I => \N__48725\
        );

    \I__11480\ : ClkMux
    port map (
            O => \N__49072\,
            I => \N__48725\
        );

    \I__11479\ : ClkMux
    port map (
            O => \N__49071\,
            I => \N__48725\
        );

    \I__11478\ : ClkMux
    port map (
            O => \N__49070\,
            I => \N__48725\
        );

    \I__11477\ : ClkMux
    port map (
            O => \N__49069\,
            I => \N__48725\
        );

    \I__11476\ : ClkMux
    port map (
            O => \N__49068\,
            I => \N__48725\
        );

    \I__11475\ : ClkMux
    port map (
            O => \N__49067\,
            I => \N__48725\
        );

    \I__11474\ : ClkMux
    port map (
            O => \N__49066\,
            I => \N__48725\
        );

    \I__11473\ : ClkMux
    port map (
            O => \N__49065\,
            I => \N__48725\
        );

    \I__11472\ : ClkMux
    port map (
            O => \N__49064\,
            I => \N__48725\
        );

    \I__11471\ : ClkMux
    port map (
            O => \N__49063\,
            I => \N__48725\
        );

    \I__11470\ : ClkMux
    port map (
            O => \N__49062\,
            I => \N__48725\
        );

    \I__11469\ : ClkMux
    port map (
            O => \N__49061\,
            I => \N__48725\
        );

    \I__11468\ : ClkMux
    port map (
            O => \N__49060\,
            I => \N__48725\
        );

    \I__11467\ : ClkMux
    port map (
            O => \N__49059\,
            I => \N__48725\
        );

    \I__11466\ : ClkMux
    port map (
            O => \N__49058\,
            I => \N__48725\
        );

    \I__11465\ : ClkMux
    port map (
            O => \N__49057\,
            I => \N__48725\
        );

    \I__11464\ : ClkMux
    port map (
            O => \N__49056\,
            I => \N__48725\
        );

    \I__11463\ : ClkMux
    port map (
            O => \N__49055\,
            I => \N__48725\
        );

    \I__11462\ : ClkMux
    port map (
            O => \N__49054\,
            I => \N__48725\
        );

    \I__11461\ : ClkMux
    port map (
            O => \N__49053\,
            I => \N__48725\
        );

    \I__11460\ : ClkMux
    port map (
            O => \N__49052\,
            I => \N__48725\
        );

    \I__11459\ : ClkMux
    port map (
            O => \N__49051\,
            I => \N__48725\
        );

    \I__11458\ : ClkMux
    port map (
            O => \N__49050\,
            I => \N__48725\
        );

    \I__11457\ : ClkMux
    port map (
            O => \N__49049\,
            I => \N__48725\
        );

    \I__11456\ : ClkMux
    port map (
            O => \N__49048\,
            I => \N__48725\
        );

    \I__11455\ : ClkMux
    port map (
            O => \N__49047\,
            I => \N__48725\
        );

    \I__11454\ : ClkMux
    port map (
            O => \N__49046\,
            I => \N__48725\
        );

    \I__11453\ : ClkMux
    port map (
            O => \N__49045\,
            I => \N__48725\
        );

    \I__11452\ : ClkMux
    port map (
            O => \N__49044\,
            I => \N__48725\
        );

    \I__11451\ : ClkMux
    port map (
            O => \N__49043\,
            I => \N__48725\
        );

    \I__11450\ : ClkMux
    port map (
            O => \N__49042\,
            I => \N__48725\
        );

    \I__11449\ : ClkMux
    port map (
            O => \N__49041\,
            I => \N__48725\
        );

    \I__11448\ : ClkMux
    port map (
            O => \N__49040\,
            I => \N__48725\
        );

    \I__11447\ : ClkMux
    port map (
            O => \N__49039\,
            I => \N__48725\
        );

    \I__11446\ : ClkMux
    port map (
            O => \N__49038\,
            I => \N__48725\
        );

    \I__11445\ : ClkMux
    port map (
            O => \N__49037\,
            I => \N__48725\
        );

    \I__11444\ : ClkMux
    port map (
            O => \N__49036\,
            I => \N__48725\
        );

    \I__11443\ : ClkMux
    port map (
            O => \N__49035\,
            I => \N__48725\
        );

    \I__11442\ : ClkMux
    port map (
            O => \N__49034\,
            I => \N__48725\
        );

    \I__11441\ : ClkMux
    port map (
            O => \N__49033\,
            I => \N__48725\
        );

    \I__11440\ : ClkMux
    port map (
            O => \N__49032\,
            I => \N__48725\
        );

    \I__11439\ : ClkMux
    port map (
            O => \N__49031\,
            I => \N__48725\
        );

    \I__11438\ : ClkMux
    port map (
            O => \N__49030\,
            I => \N__48725\
        );

    \I__11437\ : ClkMux
    port map (
            O => \N__49029\,
            I => \N__48725\
        );

    \I__11436\ : ClkMux
    port map (
            O => \N__49028\,
            I => \N__48725\
        );

    \I__11435\ : ClkMux
    port map (
            O => \N__49027\,
            I => \N__48725\
        );

    \I__11434\ : ClkMux
    port map (
            O => \N__49026\,
            I => \N__48725\
        );

    \I__11433\ : ClkMux
    port map (
            O => \N__49025\,
            I => \N__48725\
        );

    \I__11432\ : ClkMux
    port map (
            O => \N__49024\,
            I => \N__48725\
        );

    \I__11431\ : ClkMux
    port map (
            O => \N__49023\,
            I => \N__48725\
        );

    \I__11430\ : ClkMux
    port map (
            O => \N__49022\,
            I => \N__48725\
        );

    \I__11429\ : ClkMux
    port map (
            O => \N__49021\,
            I => \N__48725\
        );

    \I__11428\ : ClkMux
    port map (
            O => \N__49020\,
            I => \N__48725\
        );

    \I__11427\ : ClkMux
    port map (
            O => \N__49019\,
            I => \N__48725\
        );

    \I__11426\ : ClkMux
    port map (
            O => \N__49018\,
            I => \N__48725\
        );

    \I__11425\ : ClkMux
    port map (
            O => \N__49017\,
            I => \N__48725\
        );

    \I__11424\ : ClkMux
    port map (
            O => \N__49016\,
            I => \N__48725\
        );

    \I__11423\ : ClkMux
    port map (
            O => \N__49015\,
            I => \N__48725\
        );

    \I__11422\ : ClkMux
    port map (
            O => \N__49014\,
            I => \N__48725\
        );

    \I__11421\ : ClkMux
    port map (
            O => \N__49013\,
            I => \N__48725\
        );

    \I__11420\ : ClkMux
    port map (
            O => \N__49012\,
            I => \N__48725\
        );

    \I__11419\ : ClkMux
    port map (
            O => \N__49011\,
            I => \N__48725\
        );

    \I__11418\ : ClkMux
    port map (
            O => \N__49010\,
            I => \N__48725\
        );

    \I__11417\ : ClkMux
    port map (
            O => \N__49009\,
            I => \N__48725\
        );

    \I__11416\ : ClkMux
    port map (
            O => \N__49008\,
            I => \N__48725\
        );

    \I__11415\ : GlobalMux
    port map (
            O => \N__48725\,
            I => clk_100mhz_0
        );

    \I__11414\ : CEMux
    port map (
            O => \N__48722\,
            I => \N__48689\
        );

    \I__11413\ : CEMux
    port map (
            O => \N__48721\,
            I => \N__48689\
        );

    \I__11412\ : CEMux
    port map (
            O => \N__48720\,
            I => \N__48689\
        );

    \I__11411\ : CEMux
    port map (
            O => \N__48719\,
            I => \N__48689\
        );

    \I__11410\ : CEMux
    port map (
            O => \N__48718\,
            I => \N__48689\
        );

    \I__11409\ : CEMux
    port map (
            O => \N__48717\,
            I => \N__48689\
        );

    \I__11408\ : CEMux
    port map (
            O => \N__48716\,
            I => \N__48689\
        );

    \I__11407\ : CEMux
    port map (
            O => \N__48715\,
            I => \N__48689\
        );

    \I__11406\ : CEMux
    port map (
            O => \N__48714\,
            I => \N__48689\
        );

    \I__11405\ : CEMux
    port map (
            O => \N__48713\,
            I => \N__48689\
        );

    \I__11404\ : CEMux
    port map (
            O => \N__48712\,
            I => \N__48689\
        );

    \I__11403\ : GlobalMux
    port map (
            O => \N__48689\,
            I => \N__48686\
        );

    \I__11402\ : gio2CtrlBuf
    port map (
            O => \N__48686\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__11401\ : InMux
    port map (
            O => \N__48683\,
            I => \N__48677\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48682\,
            I => \N__48674\
        );

    \I__11399\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48671\
        );

    \I__11398\ : InMux
    port map (
            O => \N__48680\,
            I => \N__48668\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48677\,
            I => \N__48665\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__48674\,
            I => \N__48662\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48671\,
            I => \N__48659\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__48668\,
            I => \N__48560\
        );

    \I__11393\ : Glb2LocalMux
    port map (
            O => \N__48665\,
            I => \N__48227\
        );

    \I__11392\ : Glb2LocalMux
    port map (
            O => \N__48662\,
            I => \N__48227\
        );

    \I__11391\ : Glb2LocalMux
    port map (
            O => \N__48659\,
            I => \N__48227\
        );

    \I__11390\ : SRMux
    port map (
            O => \N__48658\,
            I => \N__48227\
        );

    \I__11389\ : SRMux
    port map (
            O => \N__48657\,
            I => \N__48227\
        );

    \I__11388\ : SRMux
    port map (
            O => \N__48656\,
            I => \N__48227\
        );

    \I__11387\ : SRMux
    port map (
            O => \N__48655\,
            I => \N__48227\
        );

    \I__11386\ : SRMux
    port map (
            O => \N__48654\,
            I => \N__48227\
        );

    \I__11385\ : SRMux
    port map (
            O => \N__48653\,
            I => \N__48227\
        );

    \I__11384\ : SRMux
    port map (
            O => \N__48652\,
            I => \N__48227\
        );

    \I__11383\ : SRMux
    port map (
            O => \N__48651\,
            I => \N__48227\
        );

    \I__11382\ : SRMux
    port map (
            O => \N__48650\,
            I => \N__48227\
        );

    \I__11381\ : SRMux
    port map (
            O => \N__48649\,
            I => \N__48227\
        );

    \I__11380\ : SRMux
    port map (
            O => \N__48648\,
            I => \N__48227\
        );

    \I__11379\ : SRMux
    port map (
            O => \N__48647\,
            I => \N__48227\
        );

    \I__11378\ : SRMux
    port map (
            O => \N__48646\,
            I => \N__48227\
        );

    \I__11377\ : SRMux
    port map (
            O => \N__48645\,
            I => \N__48227\
        );

    \I__11376\ : SRMux
    port map (
            O => \N__48644\,
            I => \N__48227\
        );

    \I__11375\ : SRMux
    port map (
            O => \N__48643\,
            I => \N__48227\
        );

    \I__11374\ : SRMux
    port map (
            O => \N__48642\,
            I => \N__48227\
        );

    \I__11373\ : SRMux
    port map (
            O => \N__48641\,
            I => \N__48227\
        );

    \I__11372\ : SRMux
    port map (
            O => \N__48640\,
            I => \N__48227\
        );

    \I__11371\ : SRMux
    port map (
            O => \N__48639\,
            I => \N__48227\
        );

    \I__11370\ : SRMux
    port map (
            O => \N__48638\,
            I => \N__48227\
        );

    \I__11369\ : SRMux
    port map (
            O => \N__48637\,
            I => \N__48227\
        );

    \I__11368\ : SRMux
    port map (
            O => \N__48636\,
            I => \N__48227\
        );

    \I__11367\ : SRMux
    port map (
            O => \N__48635\,
            I => \N__48227\
        );

    \I__11366\ : SRMux
    port map (
            O => \N__48634\,
            I => \N__48227\
        );

    \I__11365\ : SRMux
    port map (
            O => \N__48633\,
            I => \N__48227\
        );

    \I__11364\ : SRMux
    port map (
            O => \N__48632\,
            I => \N__48227\
        );

    \I__11363\ : SRMux
    port map (
            O => \N__48631\,
            I => \N__48227\
        );

    \I__11362\ : SRMux
    port map (
            O => \N__48630\,
            I => \N__48227\
        );

    \I__11361\ : SRMux
    port map (
            O => \N__48629\,
            I => \N__48227\
        );

    \I__11360\ : SRMux
    port map (
            O => \N__48628\,
            I => \N__48227\
        );

    \I__11359\ : SRMux
    port map (
            O => \N__48627\,
            I => \N__48227\
        );

    \I__11358\ : SRMux
    port map (
            O => \N__48626\,
            I => \N__48227\
        );

    \I__11357\ : SRMux
    port map (
            O => \N__48625\,
            I => \N__48227\
        );

    \I__11356\ : SRMux
    port map (
            O => \N__48624\,
            I => \N__48227\
        );

    \I__11355\ : SRMux
    port map (
            O => \N__48623\,
            I => \N__48227\
        );

    \I__11354\ : SRMux
    port map (
            O => \N__48622\,
            I => \N__48227\
        );

    \I__11353\ : SRMux
    port map (
            O => \N__48621\,
            I => \N__48227\
        );

    \I__11352\ : SRMux
    port map (
            O => \N__48620\,
            I => \N__48227\
        );

    \I__11351\ : SRMux
    port map (
            O => \N__48619\,
            I => \N__48227\
        );

    \I__11350\ : SRMux
    port map (
            O => \N__48618\,
            I => \N__48227\
        );

    \I__11349\ : SRMux
    port map (
            O => \N__48617\,
            I => \N__48227\
        );

    \I__11348\ : SRMux
    port map (
            O => \N__48616\,
            I => \N__48227\
        );

    \I__11347\ : SRMux
    port map (
            O => \N__48615\,
            I => \N__48227\
        );

    \I__11346\ : SRMux
    port map (
            O => \N__48614\,
            I => \N__48227\
        );

    \I__11345\ : SRMux
    port map (
            O => \N__48613\,
            I => \N__48227\
        );

    \I__11344\ : SRMux
    port map (
            O => \N__48612\,
            I => \N__48227\
        );

    \I__11343\ : SRMux
    port map (
            O => \N__48611\,
            I => \N__48227\
        );

    \I__11342\ : SRMux
    port map (
            O => \N__48610\,
            I => \N__48227\
        );

    \I__11341\ : SRMux
    port map (
            O => \N__48609\,
            I => \N__48227\
        );

    \I__11340\ : SRMux
    port map (
            O => \N__48608\,
            I => \N__48227\
        );

    \I__11339\ : SRMux
    port map (
            O => \N__48607\,
            I => \N__48227\
        );

    \I__11338\ : SRMux
    port map (
            O => \N__48606\,
            I => \N__48227\
        );

    \I__11337\ : SRMux
    port map (
            O => \N__48605\,
            I => \N__48227\
        );

    \I__11336\ : SRMux
    port map (
            O => \N__48604\,
            I => \N__48227\
        );

    \I__11335\ : SRMux
    port map (
            O => \N__48603\,
            I => \N__48227\
        );

    \I__11334\ : SRMux
    port map (
            O => \N__48602\,
            I => \N__48227\
        );

    \I__11333\ : SRMux
    port map (
            O => \N__48601\,
            I => \N__48227\
        );

    \I__11332\ : SRMux
    port map (
            O => \N__48600\,
            I => \N__48227\
        );

    \I__11331\ : SRMux
    port map (
            O => \N__48599\,
            I => \N__48227\
        );

    \I__11330\ : SRMux
    port map (
            O => \N__48598\,
            I => \N__48227\
        );

    \I__11329\ : SRMux
    port map (
            O => \N__48597\,
            I => \N__48227\
        );

    \I__11328\ : SRMux
    port map (
            O => \N__48596\,
            I => \N__48227\
        );

    \I__11327\ : SRMux
    port map (
            O => \N__48595\,
            I => \N__48227\
        );

    \I__11326\ : SRMux
    port map (
            O => \N__48594\,
            I => \N__48227\
        );

    \I__11325\ : SRMux
    port map (
            O => \N__48593\,
            I => \N__48227\
        );

    \I__11324\ : SRMux
    port map (
            O => \N__48592\,
            I => \N__48227\
        );

    \I__11323\ : SRMux
    port map (
            O => \N__48591\,
            I => \N__48227\
        );

    \I__11322\ : SRMux
    port map (
            O => \N__48590\,
            I => \N__48227\
        );

    \I__11321\ : SRMux
    port map (
            O => \N__48589\,
            I => \N__48227\
        );

    \I__11320\ : SRMux
    port map (
            O => \N__48588\,
            I => \N__48227\
        );

    \I__11319\ : SRMux
    port map (
            O => \N__48587\,
            I => \N__48227\
        );

    \I__11318\ : SRMux
    port map (
            O => \N__48586\,
            I => \N__48227\
        );

    \I__11317\ : SRMux
    port map (
            O => \N__48585\,
            I => \N__48227\
        );

    \I__11316\ : SRMux
    port map (
            O => \N__48584\,
            I => \N__48227\
        );

    \I__11315\ : SRMux
    port map (
            O => \N__48583\,
            I => \N__48227\
        );

    \I__11314\ : SRMux
    port map (
            O => \N__48582\,
            I => \N__48227\
        );

    \I__11313\ : SRMux
    port map (
            O => \N__48581\,
            I => \N__48227\
        );

    \I__11312\ : SRMux
    port map (
            O => \N__48580\,
            I => \N__48227\
        );

    \I__11311\ : SRMux
    port map (
            O => \N__48579\,
            I => \N__48227\
        );

    \I__11310\ : SRMux
    port map (
            O => \N__48578\,
            I => \N__48227\
        );

    \I__11309\ : SRMux
    port map (
            O => \N__48577\,
            I => \N__48227\
        );

    \I__11308\ : SRMux
    port map (
            O => \N__48576\,
            I => \N__48227\
        );

    \I__11307\ : SRMux
    port map (
            O => \N__48575\,
            I => \N__48227\
        );

    \I__11306\ : SRMux
    port map (
            O => \N__48574\,
            I => \N__48227\
        );

    \I__11305\ : SRMux
    port map (
            O => \N__48573\,
            I => \N__48227\
        );

    \I__11304\ : SRMux
    port map (
            O => \N__48572\,
            I => \N__48227\
        );

    \I__11303\ : SRMux
    port map (
            O => \N__48571\,
            I => \N__48227\
        );

    \I__11302\ : SRMux
    port map (
            O => \N__48570\,
            I => \N__48227\
        );

    \I__11301\ : SRMux
    port map (
            O => \N__48569\,
            I => \N__48227\
        );

    \I__11300\ : SRMux
    port map (
            O => \N__48568\,
            I => \N__48227\
        );

    \I__11299\ : SRMux
    port map (
            O => \N__48567\,
            I => \N__48227\
        );

    \I__11298\ : SRMux
    port map (
            O => \N__48566\,
            I => \N__48227\
        );

    \I__11297\ : SRMux
    port map (
            O => \N__48565\,
            I => \N__48227\
        );

    \I__11296\ : SRMux
    port map (
            O => \N__48564\,
            I => \N__48227\
        );

    \I__11295\ : SRMux
    port map (
            O => \N__48563\,
            I => \N__48227\
        );

    \I__11294\ : Glb2LocalMux
    port map (
            O => \N__48560\,
            I => \N__48227\
        );

    \I__11293\ : SRMux
    port map (
            O => \N__48559\,
            I => \N__48227\
        );

    \I__11292\ : SRMux
    port map (
            O => \N__48558\,
            I => \N__48227\
        );

    \I__11291\ : SRMux
    port map (
            O => \N__48557\,
            I => \N__48227\
        );

    \I__11290\ : SRMux
    port map (
            O => \N__48556\,
            I => \N__48227\
        );

    \I__11289\ : SRMux
    port map (
            O => \N__48555\,
            I => \N__48227\
        );

    \I__11288\ : SRMux
    port map (
            O => \N__48554\,
            I => \N__48227\
        );

    \I__11287\ : SRMux
    port map (
            O => \N__48553\,
            I => \N__48227\
        );

    \I__11286\ : SRMux
    port map (
            O => \N__48552\,
            I => \N__48227\
        );

    \I__11285\ : SRMux
    port map (
            O => \N__48551\,
            I => \N__48227\
        );

    \I__11284\ : SRMux
    port map (
            O => \N__48550\,
            I => \N__48227\
        );

    \I__11283\ : SRMux
    port map (
            O => \N__48549\,
            I => \N__48227\
        );

    \I__11282\ : SRMux
    port map (
            O => \N__48548\,
            I => \N__48227\
        );

    \I__11281\ : SRMux
    port map (
            O => \N__48547\,
            I => \N__48227\
        );

    \I__11280\ : SRMux
    port map (
            O => \N__48546\,
            I => \N__48227\
        );

    \I__11279\ : SRMux
    port map (
            O => \N__48545\,
            I => \N__48227\
        );

    \I__11278\ : SRMux
    port map (
            O => \N__48544\,
            I => \N__48227\
        );

    \I__11277\ : SRMux
    port map (
            O => \N__48543\,
            I => \N__48227\
        );

    \I__11276\ : SRMux
    port map (
            O => \N__48542\,
            I => \N__48227\
        );

    \I__11275\ : SRMux
    port map (
            O => \N__48541\,
            I => \N__48227\
        );

    \I__11274\ : SRMux
    port map (
            O => \N__48540\,
            I => \N__48227\
        );

    \I__11273\ : SRMux
    port map (
            O => \N__48539\,
            I => \N__48227\
        );

    \I__11272\ : SRMux
    port map (
            O => \N__48538\,
            I => \N__48227\
        );

    \I__11271\ : SRMux
    port map (
            O => \N__48537\,
            I => \N__48227\
        );

    \I__11270\ : SRMux
    port map (
            O => \N__48536\,
            I => \N__48227\
        );

    \I__11269\ : SRMux
    port map (
            O => \N__48535\,
            I => \N__48227\
        );

    \I__11268\ : SRMux
    port map (
            O => \N__48534\,
            I => \N__48227\
        );

    \I__11267\ : SRMux
    port map (
            O => \N__48533\,
            I => \N__48227\
        );

    \I__11266\ : SRMux
    port map (
            O => \N__48532\,
            I => \N__48227\
        );

    \I__11265\ : SRMux
    port map (
            O => \N__48531\,
            I => \N__48227\
        );

    \I__11264\ : SRMux
    port map (
            O => \N__48530\,
            I => \N__48227\
        );

    \I__11263\ : SRMux
    port map (
            O => \N__48529\,
            I => \N__48227\
        );

    \I__11262\ : SRMux
    port map (
            O => \N__48528\,
            I => \N__48227\
        );

    \I__11261\ : SRMux
    port map (
            O => \N__48527\,
            I => \N__48227\
        );

    \I__11260\ : SRMux
    port map (
            O => \N__48526\,
            I => \N__48227\
        );

    \I__11259\ : SRMux
    port map (
            O => \N__48525\,
            I => \N__48227\
        );

    \I__11258\ : SRMux
    port map (
            O => \N__48524\,
            I => \N__48227\
        );

    \I__11257\ : SRMux
    port map (
            O => \N__48523\,
            I => \N__48227\
        );

    \I__11256\ : SRMux
    port map (
            O => \N__48522\,
            I => \N__48227\
        );

    \I__11255\ : SRMux
    port map (
            O => \N__48521\,
            I => \N__48227\
        );

    \I__11254\ : SRMux
    port map (
            O => \N__48520\,
            I => \N__48227\
        );

    \I__11253\ : SRMux
    port map (
            O => \N__48519\,
            I => \N__48227\
        );

    \I__11252\ : SRMux
    port map (
            O => \N__48518\,
            I => \N__48227\
        );

    \I__11251\ : SRMux
    port map (
            O => \N__48517\,
            I => \N__48227\
        );

    \I__11250\ : SRMux
    port map (
            O => \N__48516\,
            I => \N__48227\
        );

    \I__11249\ : GlobalMux
    port map (
            O => \N__48227\,
            I => \N__48224\
        );

    \I__11248\ : gio2CtrlBuf
    port map (
            O => \N__48224\,
            I => red_c_g
        );

    \I__11247\ : InMux
    port map (
            O => \N__48221\,
            I => \N__48218\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__48218\,
            I => \N__48215\
        );

    \I__11245\ : Span4Mux_v
    port map (
            O => \N__48215\,
            I => \N__48211\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48208\
        );

    \I__11243\ : Odrv4
    port map (
            O => \N__48211\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__48208\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__11241\ : CascadeMux
    port map (
            O => \N__48203\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48200\,
            I => \N__48194\
        );

    \I__11239\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48194\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48194\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48188\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48188\,
            I => \N__48185\
        );

    \I__11235\ : Span4Mux_v
    port map (
            O => \N__48185\,
            I => \N__48182\
        );

    \I__11234\ : Odrv4
    port map (
            O => \N__48182\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48179\,
            I => \N__48173\
        );

    \I__11232\ : InMux
    port map (
            O => \N__48178\,
            I => \N__48173\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48173\,
            I => \N__48169\
        );

    \I__11230\ : InMux
    port map (
            O => \N__48172\,
            I => \N__48165\
        );

    \I__11229\ : Span4Mux_v
    port map (
            O => \N__48169\,
            I => \N__48162\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48168\,
            I => \N__48159\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__48165\,
            I => \N__48152\
        );

    \I__11226\ : Span4Mux_v
    port map (
            O => \N__48162\,
            I => \N__48152\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__48159\,
            I => \N__48152\
        );

    \I__11224\ : Odrv4
    port map (
            O => \N__48152\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__11223\ : InMux
    port map (
            O => \N__48149\,
            I => \N__48144\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48148\,
            I => \N__48140\
        );

    \I__11221\ : InMux
    port map (
            O => \N__48147\,
            I => \N__48137\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48144\,
            I => \N__48134\
        );

    \I__11219\ : InMux
    port map (
            O => \N__48143\,
            I => \N__48131\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48126\
        );

    \I__11217\ : LocalMux
    port map (
            O => \N__48137\,
            I => \N__48126\
        );

    \I__11216\ : Span4Mux_h
    port map (
            O => \N__48134\,
            I => \N__48121\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__48131\,
            I => \N__48121\
        );

    \I__11214\ : Span4Mux_v
    port map (
            O => \N__48126\,
            I => \N__48118\
        );

    \I__11213\ : Odrv4
    port map (
            O => \N__48121\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__11212\ : Odrv4
    port map (
            O => \N__48118\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__11211\ : CascadeMux
    port map (
            O => \N__48113\,
            I => \N__48108\
        );

    \I__11210\ : InMux
    port map (
            O => \N__48112\,
            I => \N__48104\
        );

    \I__11209\ : InMux
    port map (
            O => \N__48111\,
            I => \N__48101\
        );

    \I__11208\ : InMux
    port map (
            O => \N__48108\,
            I => \N__48098\
        );

    \I__11207\ : InMux
    port map (
            O => \N__48107\,
            I => \N__48095\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48104\,
            I => \N__48092\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__48087\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__48098\,
            I => \N__48087\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__48095\,
            I => \N__48084\
        );

    \I__11202\ : Span4Mux_v
    port map (
            O => \N__48092\,
            I => \N__48079\
        );

    \I__11201\ : Span4Mux_v
    port map (
            O => \N__48087\,
            I => \N__48079\
        );

    \I__11200\ : Odrv12
    port map (
            O => \N__48084\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__11199\ : Odrv4
    port map (
            O => \N__48079\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__11198\ : InMux
    port map (
            O => \N__48074\,
            I => \N__48067\
        );

    \I__11197\ : InMux
    port map (
            O => \N__48073\,
            I => \N__48067\
        );

    \I__11196\ : InMux
    port map (
            O => \N__48072\,
            I => \N__48063\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__48067\,
            I => \N__48060\
        );

    \I__11194\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48057\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__48063\,
            I => \N__48054\
        );

    \I__11192\ : Span4Mux_v
    port map (
            O => \N__48060\,
            I => \N__48049\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__48057\,
            I => \N__48049\
        );

    \I__11190\ : Odrv4
    port map (
            O => \N__48054\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__11189\ : Odrv4
    port map (
            O => \N__48049\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__11188\ : InMux
    port map (
            O => \N__48044\,
            I => \N__48041\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__48041\,
            I => \N__48038\
        );

    \I__11186\ : Odrv4
    port map (
            O => \N__48038\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__11185\ : InMux
    port map (
            O => \N__48035\,
            I => \N__48032\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__48032\,
            I => \N__48029\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__48029\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__11182\ : CascadeMux
    port map (
            O => \N__48026\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\
        );

    \I__11181\ : CascadeMux
    port map (
            O => \N__48023\,
            I => \N__48020\
        );

    \I__11180\ : InMux
    port map (
            O => \N__48020\,
            I => \N__48017\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__48017\,
            I => \N__48014\
        );

    \I__11178\ : Span4Mux_h
    port map (
            O => \N__48014\,
            I => \N__48011\
        );

    \I__11177\ : Span4Mux_h
    port map (
            O => \N__48011\,
            I => \N__48008\
        );

    \I__11176\ : Odrv4
    port map (
            O => \N__48008\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__11175\ : InMux
    port map (
            O => \N__48005\,
            I => \N__48000\
        );

    \I__11174\ : InMux
    port map (
            O => \N__48004\,
            I => \N__47995\
        );

    \I__11173\ : InMux
    port map (
            O => \N__48003\,
            I => \N__47995\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__48000\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__47995\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47990\,
            I => \N__47985\
        );

    \I__11169\ : InMux
    port map (
            O => \N__47989\,
            I => \N__47980\
        );

    \I__11168\ : InMux
    port map (
            O => \N__47988\,
            I => \N__47980\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__47985\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__47980\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__11165\ : CascadeMux
    port map (
            O => \N__47975\,
            I => \N__47972\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47972\,
            I => \N__47969\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__47969\,
            I => \N__47966\
        );

    \I__11162\ : Span4Mux_v
    port map (
            O => \N__47966\,
            I => \N__47963\
        );

    \I__11161\ : Odrv4
    port map (
            O => \N__47963\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47960\,
            I => \N__47955\
        );

    \I__11159\ : InMux
    port map (
            O => \N__47959\,
            I => \N__47952\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47958\,
            I => \N__47949\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__47955\,
            I => \N__47945\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__47952\,
            I => \N__47942\
        );

    \I__11155\ : LocalMux
    port map (
            O => \N__47949\,
            I => \N__47939\
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__47948\,
            I => \N__47936\
        );

    \I__11153\ : Span4Mux_h
    port map (
            O => \N__47945\,
            I => \N__47931\
        );

    \I__11152\ : Span4Mux_h
    port map (
            O => \N__47942\,
            I => \N__47931\
        );

    \I__11151\ : Span4Mux_h
    port map (
            O => \N__47939\,
            I => \N__47928\
        );

    \I__11150\ : InMux
    port map (
            O => \N__47936\,
            I => \N__47925\
        );

    \I__11149\ : Odrv4
    port map (
            O => \N__47931\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__11148\ : Odrv4
    port map (
            O => \N__47928\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__47925\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__11146\ : InMux
    port map (
            O => \N__47918\,
            I => \N__47915\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__47915\,
            I => \N__47910\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47914\,
            I => \N__47907\
        );

    \I__11143\ : InMux
    port map (
            O => \N__47913\,
            I => \N__47904\
        );

    \I__11142\ : Span4Mux_h
    port map (
            O => \N__47910\,
            I => \N__47901\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__47907\,
            I => \N__47898\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__47904\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__11139\ : Odrv4
    port map (
            O => \N__47901\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__11138\ : Odrv4
    port map (
            O => \N__47898\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__11137\ : InMux
    port map (
            O => \N__47891\,
            I => \N__47887\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47882\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__47887\,
            I => \N__47879\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47886\,
            I => \N__47876\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47873\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47870\
        );

    \I__11131\ : Span4Mux_h
    port map (
            O => \N__47879\,
            I => \N__47867\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47876\,
            I => \N__47864\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__47873\,
            I => \N__47861\
        );

    \I__11128\ : Odrv12
    port map (
            O => \N__47870\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__11127\ : Odrv4
    port map (
            O => \N__47867\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__11126\ : Odrv4
    port map (
            O => \N__47864\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__11125\ : Odrv4
    port map (
            O => \N__47861\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__11124\ : InMux
    port map (
            O => \N__47852\,
            I => \N__47845\
        );

    \I__11123\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47845\
        );

    \I__11122\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47841\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__47845\,
            I => \N__47838\
        );

    \I__11120\ : InMux
    port map (
            O => \N__47844\,
            I => \N__47835\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__47841\,
            I => \N__47832\
        );

    \I__11118\ : Span4Mux_h
    port map (
            O => \N__47838\,
            I => \N__47829\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__47835\,
            I => \N__47826\
        );

    \I__11116\ : Span4Mux_h
    port map (
            O => \N__47832\,
            I => \N__47823\
        );

    \I__11115\ : Span4Mux_v
    port map (
            O => \N__47829\,
            I => \N__47820\
        );

    \I__11114\ : Span4Mux_h
    port map (
            O => \N__47826\,
            I => \N__47817\
        );

    \I__11113\ : Odrv4
    port map (
            O => \N__47823\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__11112\ : Odrv4
    port map (
            O => \N__47820\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__11111\ : Odrv4
    port map (
            O => \N__47817\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47805\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47809\,
            I => \N__47802\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47808\,
            I => \N__47798\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47805\,
            I => \N__47793\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47802\,
            I => \N__47793\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47801\,
            I => \N__47790\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47798\,
            I => \N__47787\
        );

    \I__11103\ : Span4Mux_v
    port map (
            O => \N__47793\,
            I => \N__47784\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__47790\,
            I => \N__47781\
        );

    \I__11101\ : Odrv4
    port map (
            O => \N__47787\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__11100\ : Odrv4
    port map (
            O => \N__47784\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__11099\ : Odrv4
    port map (
            O => \N__47781\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47771\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__47771\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47765\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__47765\,
            I => \N__47761\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47764\,
            I => \N__47758\
        );

    \I__11093\ : Span4Mux_h
    port map (
            O => \N__47761\,
            I => \N__47753\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__47758\,
            I => \N__47750\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47745\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47756\,
            I => \N__47745\
        );

    \I__11089\ : Odrv4
    port map (
            O => \N__47753\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11088\ : Odrv4
    port map (
            O => \N__47750\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__47745\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47738\,
            I => \N__47735\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47735\,
            I => \N__47732\
        );

    \I__11084\ : Span4Mux_h
    port map (
            O => \N__47732\,
            I => \N__47729\
        );

    \I__11083\ : Odrv4
    port map (
            O => \N__47729\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__11082\ : CascadeMux
    port map (
            O => \N__47726\,
            I => \N__47723\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47717\
        );

    \I__11080\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47717\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47717\,
            I => \N__47714\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__47714\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47708\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__47708\,
            I => \N__47704\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47700\
        );

    \I__11074\ : Span12Mux_v
    port map (
            O => \N__47704\,
            I => \N__47697\
        );

    \I__11073\ : InMux
    port map (
            O => \N__47703\,
            I => \N__47694\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__47700\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__11071\ : Odrv12
    port map (
            O => \N__47697\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__47694\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47683\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47680\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__47683\,
            I => \N__47675\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47680\,
            I => \N__47672\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47679\,
            I => \N__47669\
        );

    \I__11064\ : CascadeMux
    port map (
            O => \N__47678\,
            I => \N__47666\
        );

    \I__11063\ : Span4Mux_h
    port map (
            O => \N__47675\,
            I => \N__47663\
        );

    \I__11062\ : Span4Mux_v
    port map (
            O => \N__47672\,
            I => \N__47658\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47658\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47666\,
            I => \N__47655\
        );

    \I__11059\ : Odrv4
    port map (
            O => \N__47663\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__11058\ : Odrv4
    port map (
            O => \N__47658\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47655\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__11056\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47642\
        );

    \I__11055\ : InMux
    port map (
            O => \N__47647\,
            I => \N__47642\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__47642\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__11053\ : InMux
    port map (
            O => \N__47639\,
            I => \N__47636\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__47636\,
            I => \N__47632\
        );

    \I__11051\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47628\
        );

    \I__11050\ : Span4Mux_v
    port map (
            O => \N__47632\,
            I => \N__47625\
        );

    \I__11049\ : InMux
    port map (
            O => \N__47631\,
            I => \N__47622\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47628\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__47625\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__47622\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__11045\ : CascadeMux
    port map (
            O => \N__47615\,
            I => \N__47612\
        );

    \I__11044\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47609\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__47609\,
            I => \N__47606\
        );

    \I__11042\ : Odrv4
    port map (
            O => \N__47606\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__11041\ : InMux
    port map (
            O => \N__47603\,
            I => \N__47600\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47600\,
            I => \N__47596\
        );

    \I__11039\ : InMux
    port map (
            O => \N__47599\,
            I => \N__47592\
        );

    \I__11038\ : Span12Mux_h
    port map (
            O => \N__47596\,
            I => \N__47589\
        );

    \I__11037\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47586\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47592\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__11035\ : Odrv12
    port map (
            O => \N__47589\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__47586\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47579\,
            I => \N__47573\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47573\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47573\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__11030\ : InMux
    port map (
            O => \N__47570\,
            I => \N__47564\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47569\,
            I => \N__47564\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__47564\,
            I => \N__47561\
        );

    \I__11027\ : Odrv12
    port map (
            O => \N__47561\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__11026\ : CascadeMux
    port map (
            O => \N__47558\,
            I => \N__47555\
        );

    \I__11025\ : InMux
    port map (
            O => \N__47555\,
            I => \N__47552\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__47552\,
            I => \N__47549\
        );

    \I__11023\ : Span4Mux_h
    port map (
            O => \N__47549\,
            I => \N__47546\
        );

    \I__11022\ : Odrv4
    port map (
            O => \N__47546\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__11021\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47538\
        );

    \I__11020\ : InMux
    port map (
            O => \N__47542\,
            I => \N__47533\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47533\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__47538\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__47533\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__11016\ : CascadeMux
    port map (
            O => \N__47528\,
            I => \N__47524\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47527\,
            I => \N__47520\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47524\,
            I => \N__47515\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47523\,
            I => \N__47515\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__47520\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__47515\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__11010\ : InMux
    port map (
            O => \N__47510\,
            I => \N__47507\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__47507\,
            I => \N__47504\
        );

    \I__11008\ : Odrv4
    port map (
            O => \N__47504\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47497\
        );

    \I__11006\ : InMux
    port map (
            O => \N__47500\,
            I => \N__47494\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__47497\,
            I => \N__47490\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__47494\,
            I => \N__47487\
        );

    \I__11003\ : InMux
    port map (
            O => \N__47493\,
            I => \N__47484\
        );

    \I__11002\ : Span4Mux_h
    port map (
            O => \N__47490\,
            I => \N__47479\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__47487\,
            I => \N__47479\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__47484\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__10999\ : Odrv4
    port map (
            O => \N__47479\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__10998\ : CascadeMux
    port map (
            O => \N__47474\,
            I => \N__47471\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47465\
        );

    \I__10996\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47465\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__47465\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__10994\ : CascadeMux
    port map (
            O => \N__47462\,
            I => \N__47459\
        );

    \I__10993\ : InMux
    port map (
            O => \N__47459\,
            I => \N__47456\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__47456\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47453\,
            I => \N__47449\
        );

    \I__10990\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47446\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47449\,
            I => \N__47440\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__47446\,
            I => \N__47440\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47445\,
            I => \N__47437\
        );

    \I__10986\ : Span4Mux_h
    port map (
            O => \N__47440\,
            I => \N__47434\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47437\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__47434\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__47429\,
            I => \N__47426\
        );

    \I__10982\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47422\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47425\,
            I => \N__47419\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__47422\,
            I => \N__47413\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__47419\,
            I => \N__47413\
        );

    \I__10978\ : InMux
    port map (
            O => \N__47418\,
            I => \N__47410\
        );

    \I__10977\ : Span4Mux_h
    port map (
            O => \N__47413\,
            I => \N__47407\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__47410\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10975\ : Odrv4
    port map (
            O => \N__47407\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10974\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47399\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__47399\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47396\,
            I => \N__47393\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__47393\,
            I => \N__47389\
        );

    \I__10970\ : InMux
    port map (
            O => \N__47392\,
            I => \N__47386\
        );

    \I__10969\ : Odrv12
    port map (
            O => \N__47389\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__47386\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__10967\ : CascadeMux
    port map (
            O => \N__47381\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\
        );

    \I__10966\ : InMux
    port map (
            O => \N__47378\,
            I => \N__47373\
        );

    \I__10965\ : InMux
    port map (
            O => \N__47377\,
            I => \N__47368\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47376\,
            I => \N__47368\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__47373\,
            I => \N__47365\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47362\
        );

    \I__10961\ : Span4Mux_h
    port map (
            O => \N__47365\,
            I => \N__47357\
        );

    \I__10960\ : Span4Mux_h
    port map (
            O => \N__47362\,
            I => \N__47357\
        );

    \I__10959\ : Span4Mux_v
    port map (
            O => \N__47357\,
            I => \N__47353\
        );

    \I__10958\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47350\
        );

    \I__10957\ : Odrv4
    port map (
            O => \N__47353\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__47350\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10955\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47339\
        );

    \I__10954\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47339\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__47339\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__10952\ : CascadeMux
    port map (
            O => \N__47336\,
            I => \N__47333\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47330\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__47330\,
            I => \N__47327\
        );

    \I__10949\ : Span4Mux_h
    port map (
            O => \N__47327\,
            I => \N__47324\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__47324\,
            I => \N__47321\
        );

    \I__10947\ : Odrv4
    port map (
            O => \N__47321\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47318\,
            I => \N__47315\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__47315\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__10944\ : InMux
    port map (
            O => \N__47312\,
            I => \N__47305\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47305\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47310\,
            I => \N__47302\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47305\,
            I => \N__47299\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__47302\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__10939\ : Odrv4
    port map (
            O => \N__47299\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__47294\,
            I => \N__47290\
        );

    \I__10937\ : CascadeMux
    port map (
            O => \N__47293\,
            I => \N__47287\
        );

    \I__10936\ : InMux
    port map (
            O => \N__47290\,
            I => \N__47281\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47287\,
            I => \N__47281\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47286\,
            I => \N__47278\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47281\,
            I => \N__47275\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__47278\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__10931\ : Odrv4
    port map (
            O => \N__47275\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__10930\ : CascadeMux
    port map (
            O => \N__47270\,
            I => \N__47267\
        );

    \I__10929\ : InMux
    port map (
            O => \N__47267\,
            I => \N__47264\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__47264\,
            I => \N__47261\
        );

    \I__10927\ : Odrv4
    port map (
            O => \N__47261\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__10926\ : InMux
    port map (
            O => \N__47258\,
            I => \N__47255\
        );

    \I__10925\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47251\
        );

    \I__10924\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47247\
        );

    \I__10923\ : Span4Mux_h
    port map (
            O => \N__47251\,
            I => \N__47244\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47250\,
            I => \N__47241\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__47247\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10920\ : Odrv4
    port map (
            O => \N__47244\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__47241\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10918\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47231\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__47231\,
            I => \N__47228\
        );

    \I__10916\ : Span4Mux_h
    port map (
            O => \N__47228\,
            I => \N__47222\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47219\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47214\
        );

    \I__10913\ : InMux
    port map (
            O => \N__47225\,
            I => \N__47214\
        );

    \I__10912\ : Odrv4
    port map (
            O => \N__47222\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__47219\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__47214\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10909\ : InMux
    port map (
            O => \N__47207\,
            I => \N__47204\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__47204\,
            I => \N__47201\
        );

    \I__10907\ : Span4Mux_h
    port map (
            O => \N__47201\,
            I => \N__47198\
        );

    \I__10906\ : Odrv4
    port map (
            O => \N__47198\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__10905\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47192\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__47192\,
            I => \N__47187\
        );

    \I__10903\ : InMux
    port map (
            O => \N__47191\,
            I => \N__47184\
        );

    \I__10902\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47181\
        );

    \I__10901\ : Span4Mux_h
    port map (
            O => \N__47187\,
            I => \N__47178\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__47184\,
            I => \N__47175\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__47181\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__10898\ : Odrv4
    port map (
            O => \N__47178\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__47175\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__10896\ : CEMux
    port map (
            O => \N__47168\,
            I => \N__47144\
        );

    \I__10895\ : CEMux
    port map (
            O => \N__47167\,
            I => \N__47144\
        );

    \I__10894\ : CEMux
    port map (
            O => \N__47166\,
            I => \N__47144\
        );

    \I__10893\ : CEMux
    port map (
            O => \N__47165\,
            I => \N__47144\
        );

    \I__10892\ : CEMux
    port map (
            O => \N__47164\,
            I => \N__47144\
        );

    \I__10891\ : CEMux
    port map (
            O => \N__47163\,
            I => \N__47144\
        );

    \I__10890\ : CEMux
    port map (
            O => \N__47162\,
            I => \N__47144\
        );

    \I__10889\ : CEMux
    port map (
            O => \N__47161\,
            I => \N__47144\
        );

    \I__10888\ : GlobalMux
    port map (
            O => \N__47144\,
            I => \N__47141\
        );

    \I__10887\ : gio2CtrlBuf
    port map (
            O => \N__47141\,
            I => \current_shift_inst.timer_s1.N_167_i_g\
        );

    \I__10886\ : InMux
    port map (
            O => \N__47138\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__10885\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47131\
        );

    \I__10884\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47128\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__47131\,
            I => \N__47125\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__47128\,
            I => \N__47122\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__47125\,
            I => \N__47118\
        );

    \I__10880\ : Span4Mux_h
    port map (
            O => \N__47122\,
            I => \N__47115\
        );

    \I__10879\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47112\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__47118\,
            I => \N__47109\
        );

    \I__10877\ : Span4Mux_v
    port map (
            O => \N__47115\,
            I => \N__47106\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47103\
        );

    \I__10875\ : Odrv4
    port map (
            O => \N__47109\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10874\ : Odrv4
    port map (
            O => \N__47106\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10873\ : Odrv4
    port map (
            O => \N__47103\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10872\ : InMux
    port map (
            O => \N__47096\,
            I => \N__47091\
        );

    \I__10871\ : InMux
    port map (
            O => \N__47095\,
            I => \N__47087\
        );

    \I__10870\ : InMux
    port map (
            O => \N__47094\,
            I => \N__47084\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__47091\,
            I => \N__47081\
        );

    \I__10868\ : InMux
    port map (
            O => \N__47090\,
            I => \N__47078\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__47087\,
            I => \N__47075\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__47084\,
            I => \N__47072\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__47081\,
            I => \N__47069\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__47078\,
            I => \N__47066\
        );

    \I__10863\ : Span4Mux_h
    port map (
            O => \N__47075\,
            I => \N__47063\
        );

    \I__10862\ : Span4Mux_v
    port map (
            O => \N__47072\,
            I => \N__47060\
        );

    \I__10861\ : Span4Mux_v
    port map (
            O => \N__47069\,
            I => \N__47053\
        );

    \I__10860\ : Span4Mux_v
    port map (
            O => \N__47066\,
            I => \N__47053\
        );

    \I__10859\ : Span4Mux_h
    port map (
            O => \N__47063\,
            I => \N__47053\
        );

    \I__10858\ : Odrv4
    port map (
            O => \N__47060\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__10857\ : Odrv4
    port map (
            O => \N__47053\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__10856\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47045\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__47045\,
            I => \N__47042\
        );

    \I__10854\ : Span4Mux_v
    port map (
            O => \N__47042\,
            I => \N__47037\
        );

    \I__10853\ : InMux
    port map (
            O => \N__47041\,
            I => \N__47034\
        );

    \I__10852\ : InMux
    port map (
            O => \N__47040\,
            I => \N__47031\
        );

    \I__10851\ : Span4Mux_v
    port map (
            O => \N__47037\,
            I => \N__47028\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__47034\,
            I => \N__47025\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__47031\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__10848\ : Odrv4
    port map (
            O => \N__47028\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__47025\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__10846\ : InMux
    port map (
            O => \N__47018\,
            I => \N__47015\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__47015\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__10844\ : InMux
    port map (
            O => \N__47012\,
            I => \N__47009\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__47009\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__10842\ : InMux
    port map (
            O => \N__47006\,
            I => \N__47003\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__47003\,
            I => \N__47000\
        );

    \I__10840\ : Span4Mux_v
    port map (
            O => \N__47000\,
            I => \N__46997\
        );

    \I__10839\ : Span4Mux_h
    port map (
            O => \N__46997\,
            I => \N__46993\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46996\,
            I => \N__46990\
        );

    \I__10837\ : Odrv4
    port map (
            O => \N__46993\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__46990\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10835\ : CascadeMux
    port map (
            O => \N__46985\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__10834\ : InMux
    port map (
            O => \N__46982\,
            I => \N__46976\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46981\,
            I => \N__46976\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46976\,
            I => \N__46972\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46969\
        );

    \I__10830\ : Span4Mux_h
    port map (
            O => \N__46972\,
            I => \N__46966\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__46969\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10828\ : Odrv4
    port map (
            O => \N__46966\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10827\ : CascadeMux
    port map (
            O => \N__46961\,
            I => \N__46957\
        );

    \I__10826\ : CascadeMux
    port map (
            O => \N__46960\,
            I => \N__46954\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46949\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46954\,
            I => \N__46949\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__46949\,
            I => \N__46945\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46948\,
            I => \N__46942\
        );

    \I__10821\ : Span4Mux_h
    port map (
            O => \N__46945\,
            I => \N__46939\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46942\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__46939\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46928\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46933\,
            I => \N__46928\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__46928\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__10815\ : CascadeMux
    port map (
            O => \N__46925\,
            I => \N__46922\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46919\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46919\,
            I => \N__46916\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__46916\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46913\,
            I => \N__46910\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46910\,
            I => \N__46907\
        );

    \I__10809\ : Span4Mux_v
    port map (
            O => \N__46907\,
            I => \N__46903\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46900\
        );

    \I__10807\ : Odrv4
    port map (
            O => \N__46903\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46900\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10805\ : CascadeMux
    port map (
            O => \N__46895\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46889\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__46889\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__10802\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46880\
        );

    \I__10801\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46880\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__46880\,
            I => \N__46876\
        );

    \I__10799\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46873\
        );

    \I__10798\ : Span4Mux_h
    port map (
            O => \N__46876\,
            I => \N__46870\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__46873\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10796\ : Odrv4
    port map (
            O => \N__46870\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10795\ : CascadeMux
    port map (
            O => \N__46865\,
            I => \N__46862\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46862\,
            I => \N__46858\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46861\,
            I => \N__46855\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__46858\,
            I => \N__46851\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46855\,
            I => \N__46848\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46854\,
            I => \N__46845\
        );

    \I__10789\ : Span4Mux_h
    port map (
            O => \N__46851\,
            I => \N__46840\
        );

    \I__10788\ : Span4Mux_h
    port map (
            O => \N__46848\,
            I => \N__46840\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46837\
        );

    \I__10786\ : Span4Mux_v
    port map (
            O => \N__46840\,
            I => \N__46833\
        );

    \I__10785\ : Span4Mux_h
    port map (
            O => \N__46837\,
            I => \N__46830\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46836\,
            I => \N__46827\
        );

    \I__10783\ : Odrv4
    port map (
            O => \N__46833\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10782\ : Odrv4
    port map (
            O => \N__46830\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46827\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46820\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46811\
        );

    \I__10778\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46811\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46811\,
            I => \N__46807\
        );

    \I__10776\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46804\
        );

    \I__10775\ : Span4Mux_h
    port map (
            O => \N__46807\,
            I => \N__46801\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__46804\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10773\ : Odrv4
    port map (
            O => \N__46801\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10772\ : CascadeMux
    port map (
            O => \N__46796\,
            I => \N__46792\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46789\
        );

    \I__10770\ : InMux
    port map (
            O => \N__46792\,
            I => \N__46786\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__46789\,
            I => \N__46783\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46786\,
            I => \N__46779\
        );

    \I__10767\ : Span4Mux_h
    port map (
            O => \N__46783\,
            I => \N__46776\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46782\,
            I => \N__46773\
        );

    \I__10765\ : Span4Mux_h
    port map (
            O => \N__46779\,
            I => \N__46767\
        );

    \I__10764\ : Span4Mux_v
    port map (
            O => \N__46776\,
            I => \N__46767\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46764\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46761\
        );

    \I__10761\ : Odrv4
    port map (
            O => \N__46767\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10760\ : Odrv4
    port map (
            O => \N__46764\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46761\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46754\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__46751\,
            I => \N__46747\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__46750\,
            I => \N__46744\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46739\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46739\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__46739\,
            I => \N__46735\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46738\,
            I => \N__46732\
        );

    \I__10751\ : Span4Mux_h
    port map (
            O => \N__46735\,
            I => \N__46729\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46732\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10749\ : Odrv4
    port map (
            O => \N__46729\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10748\ : CascadeMux
    port map (
            O => \N__46724\,
            I => \N__46721\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46721\,
            I => \N__46717\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46720\,
            I => \N__46713\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__46717\,
            I => \N__46710\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46707\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46713\,
            I => \N__46704\
        );

    \I__10742\ : Span4Mux_v
    port map (
            O => \N__46710\,
            I => \N__46701\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46707\,
            I => \N__46698\
        );

    \I__10740\ : Span4Mux_h
    port map (
            O => \N__46704\,
            I => \N__46694\
        );

    \I__10739\ : Span4Mux_h
    port map (
            O => \N__46701\,
            I => \N__46691\
        );

    \I__10738\ : Span12Mux_v
    port map (
            O => \N__46698\,
            I => \N__46688\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46685\
        );

    \I__10736\ : Odrv4
    port map (
            O => \N__46694\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10735\ : Odrv4
    port map (
            O => \N__46691\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10734\ : Odrv12
    port map (
            O => \N__46688\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__46685\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46676\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__10731\ : CascadeMux
    port map (
            O => \N__46673\,
            I => \N__46669\
        );

    \I__10730\ : CascadeMux
    port map (
            O => \N__46672\,
            I => \N__46666\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46669\,
            I => \N__46661\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46661\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__46661\,
            I => \N__46657\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46660\,
            I => \N__46654\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__46657\,
            I => \N__46651\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__46654\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__10723\ : Odrv4
    port map (
            O => \N__46651\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46642\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46645\,
            I => \N__46638\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__46642\,
            I => \N__46635\
        );

    \I__10719\ : InMux
    port map (
            O => \N__46641\,
            I => \N__46632\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__46638\,
            I => \N__46629\
        );

    \I__10717\ : Span4Mux_v
    port map (
            O => \N__46635\,
            I => \N__46624\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46632\,
            I => \N__46624\
        );

    \I__10715\ : Span4Mux_h
    port map (
            O => \N__46629\,
            I => \N__46620\
        );

    \I__10714\ : Span4Mux_h
    port map (
            O => \N__46624\,
            I => \N__46617\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46623\,
            I => \N__46614\
        );

    \I__10712\ : Odrv4
    port map (
            O => \N__46620\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10711\ : Odrv4
    port map (
            O => \N__46617\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__46614\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46607\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__10708\ : CascadeMux
    port map (
            O => \N__46604\,
            I => \N__46601\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46601\,
            I => \N__46598\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46598\,
            I => \N__46594\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46597\,
            I => \N__46591\
        );

    \I__10704\ : Span4Mux_v
    port map (
            O => \N__46594\,
            I => \N__46585\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__46591\,
            I => \N__46585\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46582\
        );

    \I__10701\ : Span4Mux_h
    port map (
            O => \N__46585\,
            I => \N__46579\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__46582\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10699\ : Odrv4
    port map (
            O => \N__46579\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10698\ : InMux
    port map (
            O => \N__46574\,
            I => \N__46571\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46567\
        );

    \I__10696\ : CascadeMux
    port map (
            O => \N__46570\,
            I => \N__46564\
        );

    \I__10695\ : Span4Mux_h
    port map (
            O => \N__46567\,
            I => \N__46559\
        );

    \I__10694\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46554\
        );

    \I__10693\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46554\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46551\
        );

    \I__10691\ : Span4Mux_v
    port map (
            O => \N__46559\,
            I => \N__46544\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__46554\,
            I => \N__46544\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46544\
        );

    \I__10688\ : Span4Mux_h
    port map (
            O => \N__46544\,
            I => \N__46541\
        );

    \I__10687\ : Odrv4
    port map (
            O => \N__46541\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__10686\ : InMux
    port map (
            O => \N__46538\,
            I => \bfn_18_14_0_\
        );

    \I__10685\ : CascadeMux
    port map (
            O => \N__46535\,
            I => \N__46532\
        );

    \I__10684\ : InMux
    port map (
            O => \N__46532\,
            I => \N__46529\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__46529\,
            I => \N__46525\
        );

    \I__10682\ : InMux
    port map (
            O => \N__46528\,
            I => \N__46522\
        );

    \I__10681\ : Span4Mux_v
    port map (
            O => \N__46525\,
            I => \N__46516\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__46522\,
            I => \N__46516\
        );

    \I__10679\ : InMux
    port map (
            O => \N__46521\,
            I => \N__46513\
        );

    \I__10678\ : Span4Mux_h
    port map (
            O => \N__46516\,
            I => \N__46510\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__46513\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10676\ : Odrv4
    port map (
            O => \N__46510\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10675\ : CascadeMux
    port map (
            O => \N__46505\,
            I => \N__46502\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46498\
        );

    \I__10673\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46494\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46498\,
            I => \N__46491\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46497\,
            I => \N__46488\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__46494\,
            I => \N__46485\
        );

    \I__10669\ : Span4Mux_h
    port map (
            O => \N__46491\,
            I => \N__46482\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__46488\,
            I => \N__46479\
        );

    \I__10667\ : Span4Mux_h
    port map (
            O => \N__46485\,
            I => \N__46475\
        );

    \I__10666\ : Span4Mux_v
    port map (
            O => \N__46482\,
            I => \N__46472\
        );

    \I__10665\ : Span4Mux_h
    port map (
            O => \N__46479\,
            I => \N__46469\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46466\
        );

    \I__10663\ : Odrv4
    port map (
            O => \N__46475\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__10662\ : Odrv4
    port map (
            O => \N__46472\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__10661\ : Odrv4
    port map (
            O => \N__46469\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46466\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46457\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46454\,
            I => \N__46451\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__46451\,
            I => \N__46447\
        );

    \I__10656\ : InMux
    port map (
            O => \N__46450\,
            I => \N__46444\
        );

    \I__10655\ : Span4Mux_h
    port map (
            O => \N__46447\,
            I => \N__46441\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46444\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10653\ : Odrv4
    port map (
            O => \N__46441\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10652\ : CascadeMux
    port map (
            O => \N__46436\,
            I => \N__46433\
        );

    \I__10651\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46428\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46432\,
            I => \N__46425\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46431\,
            I => \N__46422\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__46428\,
            I => \N__46417\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__46425\,
            I => \N__46417\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__46422\,
            I => \N__46412\
        );

    \I__10645\ : Span4Mux_v
    port map (
            O => \N__46417\,
            I => \N__46412\
        );

    \I__10644\ : Odrv4
    port map (
            O => \N__46412\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46403\
        );

    \I__10642\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46398\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46407\,
            I => \N__46398\
        );

    \I__10640\ : InMux
    port map (
            O => \N__46406\,
            I => \N__46395\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46403\,
            I => \N__46392\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__46398\,
            I => \N__46387\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46395\,
            I => \N__46387\
        );

    \I__10636\ : Span4Mux_h
    port map (
            O => \N__46392\,
            I => \N__46384\
        );

    \I__10635\ : Span4Mux_v
    port map (
            O => \N__46387\,
            I => \N__46381\
        );

    \I__10634\ : Odrv4
    port map (
            O => \N__46384\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__46381\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__10632\ : InMux
    port map (
            O => \N__46376\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46370\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__46370\,
            I => \N__46366\
        );

    \I__10629\ : InMux
    port map (
            O => \N__46369\,
            I => \N__46363\
        );

    \I__10628\ : Span4Mux_h
    port map (
            O => \N__46366\,
            I => \N__46360\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46363\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__46360\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10625\ : CascadeMux
    port map (
            O => \N__46355\,
            I => \N__46352\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46348\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46351\,
            I => \N__46345\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__46348\,
            I => \N__46339\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46339\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46336\
        );

    \I__10619\ : Span4Mux_v
    port map (
            O => \N__46339\,
            I => \N__46333\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__46336\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10617\ : Odrv4
    port map (
            O => \N__46333\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__46328\,
            I => \N__46325\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46325\,
            I => \N__46321\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46324\,
            I => \N__46317\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__46321\,
            I => \N__46314\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46320\,
            I => \N__46311\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__46317\,
            I => \N__46308\
        );

    \I__10610\ : Span4Mux_v
    port map (
            O => \N__46314\,
            I => \N__46303\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__46311\,
            I => \N__46303\
        );

    \I__10608\ : Span4Mux_v
    port map (
            O => \N__46308\,
            I => \N__46299\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__46303\,
            I => \N__46296\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46293\
        );

    \I__10605\ : Odrv4
    port map (
            O => \N__46299\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10604\ : Odrv4
    port map (
            O => \N__46296\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__46293\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46286\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__10601\ : CascadeMux
    port map (
            O => \N__46283\,
            I => \N__46280\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46276\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46273\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__46276\,
            I => \N__46267\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__46273\,
            I => \N__46267\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46264\
        );

    \I__10595\ : Span4Mux_h
    port map (
            O => \N__46267\,
            I => \N__46261\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__46264\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10593\ : Odrv4
    port map (
            O => \N__46261\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10592\ : CascadeMux
    port map (
            O => \N__46256\,
            I => \N__46253\
        );

    \I__10591\ : InMux
    port map (
            O => \N__46253\,
            I => \N__46249\
        );

    \I__10590\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46246\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__46249\,
            I => \N__46242\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__46246\,
            I => \N__46239\
        );

    \I__10587\ : InMux
    port map (
            O => \N__46245\,
            I => \N__46236\
        );

    \I__10586\ : Span4Mux_v
    port map (
            O => \N__46242\,
            I => \N__46229\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__46239\,
            I => \N__46229\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46236\,
            I => \N__46229\
        );

    \I__10583\ : Span4Mux_h
    port map (
            O => \N__46229\,
            I => \N__46225\
        );

    \I__10582\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46222\
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__46225\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__46222\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10579\ : InMux
    port map (
            O => \N__46217\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__10578\ : InMux
    port map (
            O => \N__46214\,
            I => \N__46208\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46208\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__46208\,
            I => \N__46204\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46207\,
            I => \N__46201\
        );

    \I__10574\ : Span4Mux_h
    port map (
            O => \N__46204\,
            I => \N__46198\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__46201\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10572\ : Odrv4
    port map (
            O => \N__46198\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10571\ : CascadeMux
    port map (
            O => \N__46193\,
            I => \N__46190\
        );

    \I__10570\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46187\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__46187\,
            I => \N__46184\
        );

    \I__10568\ : Span4Mux_v
    port map (
            O => \N__46184\,
            I => \N__46180\
        );

    \I__10567\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46177\
        );

    \I__10566\ : Span4Mux_h
    port map (
            O => \N__46180\,
            I => \N__46173\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__46177\,
            I => \N__46170\
        );

    \I__10564\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46167\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__46173\,
            I => \N__46162\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__46170\,
            I => \N__46162\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__46167\,
            I => \N__46159\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__46162\,
            I => \N__46155\
        );

    \I__10559\ : Span4Mux_h
    port map (
            O => \N__46159\,
            I => \N__46152\
        );

    \I__10558\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46149\
        );

    \I__10557\ : Odrv4
    port map (
            O => \N__46155\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10556\ : Odrv4
    port map (
            O => \N__46152\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46149\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10554\ : InMux
    port map (
            O => \N__46142\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__10553\ : CascadeMux
    port map (
            O => \N__46139\,
            I => \N__46136\
        );

    \I__10552\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46132\
        );

    \I__10551\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46129\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__46132\,
            I => \N__46123\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46123\
        );

    \I__10548\ : InMux
    port map (
            O => \N__46128\,
            I => \N__46120\
        );

    \I__10547\ : Span4Mux_h
    port map (
            O => \N__46123\,
            I => \N__46117\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__46120\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__46117\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10544\ : CascadeMux
    port map (
            O => \N__46112\,
            I => \N__46108\
        );

    \I__10543\ : CascadeMux
    port map (
            O => \N__46111\,
            I => \N__46105\
        );

    \I__10542\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46102\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46105\,
            I => \N__46098\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__46102\,
            I => \N__46095\
        );

    \I__10539\ : InMux
    port map (
            O => \N__46101\,
            I => \N__46091\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__46098\,
            I => \N__46088\
        );

    \I__10537\ : Span4Mux_v
    port map (
            O => \N__46095\,
            I => \N__46085\
        );

    \I__10536\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46082\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__46091\,
            I => \N__46079\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__46088\,
            I => \N__46072\
        );

    \I__10533\ : Span4Mux_v
    port map (
            O => \N__46085\,
            I => \N__46072\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__46082\,
            I => \N__46072\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__46079\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__46072\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10529\ : InMux
    port map (
            O => \N__46067\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__46064\,
            I => \N__46060\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__46063\,
            I => \N__46057\
        );

    \I__10526\ : InMux
    port map (
            O => \N__46060\,
            I => \N__46052\
        );

    \I__10525\ : InMux
    port map (
            O => \N__46057\,
            I => \N__46052\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__46052\,
            I => \N__46048\
        );

    \I__10523\ : InMux
    port map (
            O => \N__46051\,
            I => \N__46045\
        );

    \I__10522\ : Span4Mux_h
    port map (
            O => \N__46048\,
            I => \N__46042\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__46045\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__46042\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__10519\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46032\
        );

    \I__10518\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46029\
        );

    \I__10517\ : InMux
    port map (
            O => \N__46035\,
            I => \N__46025\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__46032\,
            I => \N__46020\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__46029\,
            I => \N__46020\
        );

    \I__10514\ : InMux
    port map (
            O => \N__46028\,
            I => \N__46017\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__46025\,
            I => \N__46014\
        );

    \I__10512\ : Span4Mux_v
    port map (
            O => \N__46020\,
            I => \N__46009\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__46017\,
            I => \N__46009\
        );

    \I__10510\ : Odrv4
    port map (
            O => \N__46014\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10509\ : Odrv4
    port map (
            O => \N__46009\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10508\ : InMux
    port map (
            O => \N__46004\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__10507\ : CascadeMux
    port map (
            O => \N__46001\,
            I => \N__45998\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45995\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__45995\,
            I => \N__45991\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45988\
        );

    \I__10503\ : Span4Mux_v
    port map (
            O => \N__45991\,
            I => \N__45982\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__45988\,
            I => \N__45982\
        );

    \I__10501\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45979\
        );

    \I__10500\ : Span4Mux_h
    port map (
            O => \N__45982\,
            I => \N__45976\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__45979\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__45976\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__10497\ : CascadeMux
    port map (
            O => \N__45971\,
            I => \N__45968\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45964\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45967\,
            I => \N__45960\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45964\,
            I => \N__45957\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45963\,
            I => \N__45954\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__45960\,
            I => \N__45951\
        );

    \I__10491\ : Span4Mux_v
    port map (
            O => \N__45957\,
            I => \N__45946\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45954\,
            I => \N__45946\
        );

    \I__10489\ : Span4Mux_v
    port map (
            O => \N__45951\,
            I => \N__45942\
        );

    \I__10488\ : Span4Mux_v
    port map (
            O => \N__45946\,
            I => \N__45939\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45945\,
            I => \N__45936\
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__45942\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10485\ : Odrv4
    port map (
            O => \N__45939\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__45936\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10483\ : InMux
    port map (
            O => \N__45929\,
            I => \bfn_18_13_0_\
        );

    \I__10482\ : CascadeMux
    port map (
            O => \N__45926\,
            I => \N__45923\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45920\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45920\,
            I => \N__45916\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45919\,
            I => \N__45913\
        );

    \I__10478\ : Span4Mux_v
    port map (
            O => \N__45916\,
            I => \N__45907\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45913\,
            I => \N__45907\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45904\
        );

    \I__10475\ : Span4Mux_h
    port map (
            O => \N__45907\,
            I => \N__45901\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45904\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__10473\ : Odrv4
    port map (
            O => \N__45901\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__10472\ : CascadeMux
    port map (
            O => \N__45896\,
            I => \N__45892\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45888\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45892\,
            I => \N__45885\
        );

    \I__10469\ : CascadeMux
    port map (
            O => \N__45891\,
            I => \N__45882\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45877\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45885\,
            I => \N__45877\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45874\
        );

    \I__10465\ : Span4Mux_h
    port map (
            O => \N__45877\,
            I => \N__45870\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__45874\,
            I => \N__45867\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45864\
        );

    \I__10462\ : Odrv4
    port map (
            O => \N__45870\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__45867\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45864\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45857\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__10458\ : CascadeMux
    port map (
            O => \N__45854\,
            I => \N__45851\
        );

    \I__10457\ : InMux
    port map (
            O => \N__45851\,
            I => \N__45847\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45850\,
            I => \N__45844\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__45847\,
            I => \N__45838\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45844\,
            I => \N__45838\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45843\,
            I => \N__45835\
        );

    \I__10452\ : Span4Mux_v
    port map (
            O => \N__45838\,
            I => \N__45832\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45835\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__10450\ : Odrv4
    port map (
            O => \N__45832\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__10449\ : CascadeMux
    port map (
            O => \N__45827\,
            I => \N__45824\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45824\,
            I => \N__45820\
        );

    \I__10447\ : InMux
    port map (
            O => \N__45823\,
            I => \N__45816\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45820\,
            I => \N__45813\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45819\,
            I => \N__45810\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__45816\,
            I => \N__45807\
        );

    \I__10443\ : Span4Mux_v
    port map (
            O => \N__45813\,
            I => \N__45804\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45810\,
            I => \N__45801\
        );

    \I__10441\ : Span4Mux_v
    port map (
            O => \N__45807\,
            I => \N__45797\
        );

    \I__10440\ : Span4Mux_v
    port map (
            O => \N__45804\,
            I => \N__45794\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__45801\,
            I => \N__45791\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45800\,
            I => \N__45788\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__45797\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10436\ : Odrv4
    port map (
            O => \N__45794\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10435\ : Odrv4
    port map (
            O => \N__45791\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__45788\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45779\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__10432\ : CascadeMux
    port map (
            O => \N__45776\,
            I => \N__45773\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45773\,
            I => \N__45768\
        );

    \I__10430\ : InMux
    port map (
            O => \N__45772\,
            I => \N__45765\
        );

    \I__10429\ : InMux
    port map (
            O => \N__45771\,
            I => \N__45762\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45768\,
            I => \N__45757\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45757\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45762\,
            I => \N__45752\
        );

    \I__10425\ : Span4Mux_v
    port map (
            O => \N__45757\,
            I => \N__45752\
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__45752\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45740\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45748\,
            I => \N__45740\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45740\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__45740\,
            I => \N__45736\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45739\,
            I => \N__45733\
        );

    \I__10418\ : Odrv4
    port map (
            O => \N__45736\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__45733\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45728\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__10415\ : CascadeMux
    port map (
            O => \N__45725\,
            I => \N__45722\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45718\
        );

    \I__10413\ : InMux
    port map (
            O => \N__45721\,
            I => \N__45715\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__45718\,
            I => \N__45709\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45715\,
            I => \N__45709\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45706\
        );

    \I__10409\ : Span4Mux_h
    port map (
            O => \N__45709\,
            I => \N__45703\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__45706\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__10407\ : Odrv4
    port map (
            O => \N__45703\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__10406\ : CascadeMux
    port map (
            O => \N__45698\,
            I => \N__45695\
        );

    \I__10405\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45691\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45688\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45684\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__45688\,
            I => \N__45681\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45687\,
            I => \N__45678\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__45684\,
            I => \N__45674\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__45681\,
            I => \N__45671\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45668\
        );

    \I__10397\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45665\
        );

    \I__10396\ : Span4Mux_v
    port map (
            O => \N__45674\,
            I => \N__45662\
        );

    \I__10395\ : Span4Mux_h
    port map (
            O => \N__45671\,
            I => \N__45655\
        );

    \I__10394\ : Span4Mux_v
    port map (
            O => \N__45668\,
            I => \N__45655\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__45665\,
            I => \N__45655\
        );

    \I__10392\ : Odrv4
    port map (
            O => \N__45662\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10391\ : Odrv4
    port map (
            O => \N__45655\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10390\ : InMux
    port map (
            O => \N__45650\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__10389\ : InMux
    port map (
            O => \N__45647\,
            I => \N__45641\
        );

    \I__10388\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45641\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__45641\,
            I => \N__45637\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45640\,
            I => \N__45634\
        );

    \I__10385\ : Span4Mux_h
    port map (
            O => \N__45637\,
            I => \N__45631\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45634\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__10383\ : Odrv4
    port map (
            O => \N__45631\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45626\,
            I => \N__45623\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__45623\,
            I => \N__45617\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45622\,
            I => \N__45612\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45612\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45620\,
            I => \N__45609\
        );

    \I__10377\ : Span4Mux_h
    port map (
            O => \N__45617\,
            I => \N__45606\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45612\,
            I => \N__45603\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__45609\,
            I => \N__45600\
        );

    \I__10374\ : Span4Mux_v
    port map (
            O => \N__45606\,
            I => \N__45597\
        );

    \I__10373\ : Span4Mux_v
    port map (
            O => \N__45603\,
            I => \N__45592\
        );

    \I__10372\ : Span4Mux_h
    port map (
            O => \N__45600\,
            I => \N__45592\
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__45597\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10370\ : Odrv4
    port map (
            O => \N__45592\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45587\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45584\,
            I => \N__45578\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45578\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__45578\,
            I => \N__45574\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45571\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__45574\,
            I => \N__45568\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__45571\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__45568\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45563\,
            I => \N__45559\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__45562\,
            I => \N__45556\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45553\
        );

    \I__10358\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45550\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__45553\,
            I => \N__45545\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__45550\,
            I => \N__45542\
        );

    \I__10355\ : InMux
    port map (
            O => \N__45549\,
            I => \N__45539\
        );

    \I__10354\ : InMux
    port map (
            O => \N__45548\,
            I => \N__45536\
        );

    \I__10353\ : Span4Mux_h
    port map (
            O => \N__45545\,
            I => \N__45531\
        );

    \I__10352\ : Span4Mux_h
    port map (
            O => \N__45542\,
            I => \N__45531\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__45539\,
            I => \N__45528\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45536\,
            I => \N__45525\
        );

    \I__10349\ : Span4Mux_v
    port map (
            O => \N__45531\,
            I => \N__45522\
        );

    \I__10348\ : Sp12to4
    port map (
            O => \N__45528\,
            I => \N__45519\
        );

    \I__10347\ : Span4Mux_h
    port map (
            O => \N__45525\,
            I => \N__45516\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__45522\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10345\ : Odrv12
    port map (
            O => \N__45519\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10344\ : Odrv4
    port map (
            O => \N__45516\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45509\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__10342\ : CascadeMux
    port map (
            O => \N__45506\,
            I => \N__45502\
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__45505\,
            I => \N__45499\
        );

    \I__10340\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45494\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45499\,
            I => \N__45494\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__45494\,
            I => \N__45490\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45487\
        );

    \I__10336\ : Span4Mux_h
    port map (
            O => \N__45490\,
            I => \N__45484\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__45487\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__10334\ : Odrv4
    port map (
            O => \N__45484\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__10333\ : InMux
    port map (
            O => \N__45479\,
            I => \N__45471\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45471\
        );

    \I__10331\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45468\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45476\,
            I => \N__45465\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45462\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__45468\,
            I => \N__45459\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__45465\,
            I => \N__45454\
        );

    \I__10326\ : Span4Mux_h
    port map (
            O => \N__45462\,
            I => \N__45454\
        );

    \I__10325\ : Span12Mux_s10_v
    port map (
            O => \N__45459\,
            I => \N__45451\
        );

    \I__10324\ : Span4Mux_h
    port map (
            O => \N__45454\,
            I => \N__45448\
        );

    \I__10323\ : Odrv12
    port map (
            O => \N__45451\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10322\ : Odrv4
    port map (
            O => \N__45448\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45443\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__10320\ : CascadeMux
    port map (
            O => \N__45440\,
            I => \N__45436\
        );

    \I__10319\ : CascadeMux
    port map (
            O => \N__45439\,
            I => \N__45433\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45430\
        );

    \I__10317\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45427\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__45430\,
            I => \N__45423\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__45427\,
            I => \N__45420\
        );

    \I__10314\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45417\
        );

    \I__10313\ : Span4Mux_h
    port map (
            O => \N__45423\,
            I => \N__45414\
        );

    \I__10312\ : Span4Mux_h
    port map (
            O => \N__45420\,
            I => \N__45411\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45417\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10310\ : Odrv4
    port map (
            O => \N__45414\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__45411\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10308\ : CascadeMux
    port map (
            O => \N__45404\,
            I => \N__45400\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45397\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45400\,
            I => \N__45394\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__45397\,
            I => \N__45390\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__45394\,
            I => \N__45387\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45384\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__45390\,
            I => \N__45379\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__45387\,
            I => \N__45379\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45384\,
            I => \N__45376\
        );

    \I__10299\ : Span4Mux_h
    port map (
            O => \N__45379\,
            I => \N__45372\
        );

    \I__10298\ : Span4Mux_h
    port map (
            O => \N__45376\,
            I => \N__45369\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45375\,
            I => \N__45366\
        );

    \I__10296\ : Odrv4
    port map (
            O => \N__45372\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10295\ : Odrv4
    port map (
            O => \N__45369\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__45366\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10293\ : InMux
    port map (
            O => \N__45359\,
            I => \bfn_18_12_0_\
        );

    \I__10292\ : CascadeMux
    port map (
            O => \N__45356\,
            I => \N__45353\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45349\
        );

    \I__10290\ : InMux
    port map (
            O => \N__45352\,
            I => \N__45346\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45349\,
            I => \N__45342\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45346\,
            I => \N__45339\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45336\
        );

    \I__10286\ : Span4Mux_h
    port map (
            O => \N__45342\,
            I => \N__45333\
        );

    \I__10285\ : Span4Mux_h
    port map (
            O => \N__45339\,
            I => \N__45330\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__45336\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__45333\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10282\ : Odrv4
    port map (
            O => \N__45330\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10281\ : CascadeMux
    port map (
            O => \N__45323\,
            I => \N__45319\
        );

    \I__10280\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45316\
        );

    \I__10279\ : InMux
    port map (
            O => \N__45319\,
            I => \N__45313\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45316\,
            I => \N__45309\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__45313\,
            I => \N__45306\
        );

    \I__10276\ : InMux
    port map (
            O => \N__45312\,
            I => \N__45303\
        );

    \I__10275\ : Span4Mux_h
    port map (
            O => \N__45309\,
            I => \N__45298\
        );

    \I__10274\ : Span4Mux_h
    port map (
            O => \N__45306\,
            I => \N__45298\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__45303\,
            I => \N__45295\
        );

    \I__10272\ : Span4Mux_v
    port map (
            O => \N__45298\,
            I => \N__45291\
        );

    \I__10271\ : Span4Mux_h
    port map (
            O => \N__45295\,
            I => \N__45288\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45285\
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__45291\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10268\ : Odrv4
    port map (
            O => \N__45288\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__45285\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10266\ : InMux
    port map (
            O => \N__45278\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__10265\ : CascadeMux
    port map (
            O => \N__45275\,
            I => \N__45272\
        );

    \I__10264\ : InMux
    port map (
            O => \N__45272\,
            I => \N__45268\
        );

    \I__10263\ : InMux
    port map (
            O => \N__45271\,
            I => \N__45265\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__45268\,
            I => \N__45259\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__45265\,
            I => \N__45259\
        );

    \I__10260\ : InMux
    port map (
            O => \N__45264\,
            I => \N__45256\
        );

    \I__10259\ : Span4Mux_v
    port map (
            O => \N__45259\,
            I => \N__45253\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__45256\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__10257\ : Odrv4
    port map (
            O => \N__45253\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__10256\ : CascadeMux
    port map (
            O => \N__45248\,
            I => \N__45244\
        );

    \I__10255\ : CascadeMux
    port map (
            O => \N__45247\,
            I => \N__45241\
        );

    \I__10254\ : InMux
    port map (
            O => \N__45244\,
            I => \N__45238\
        );

    \I__10253\ : InMux
    port map (
            O => \N__45241\,
            I => \N__45235\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__45238\,
            I => \N__45232\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__45235\,
            I => \N__45228\
        );

    \I__10250\ : Span4Mux_v
    port map (
            O => \N__45232\,
            I => \N__45225\
        );

    \I__10249\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45222\
        );

    \I__10248\ : Span4Mux_v
    port map (
            O => \N__45228\,
            I => \N__45218\
        );

    \I__10247\ : Span4Mux_v
    port map (
            O => \N__45225\,
            I => \N__45215\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__45222\,
            I => \N__45212\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45209\
        );

    \I__10244\ : Odrv4
    port map (
            O => \N__45218\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10243\ : Odrv4
    port map (
            O => \N__45215\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10242\ : Odrv4
    port map (
            O => \N__45212\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__45209\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10240\ : InMux
    port map (
            O => \N__45200\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__10239\ : CascadeMux
    port map (
            O => \N__45197\,
            I => \N__45194\
        );

    \I__10238\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45190\
        );

    \I__10237\ : InMux
    port map (
            O => \N__45193\,
            I => \N__45187\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__45190\,
            I => \N__45181\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45187\,
            I => \N__45181\
        );

    \I__10234\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45178\
        );

    \I__10233\ : Span4Mux_v
    port map (
            O => \N__45181\,
            I => \N__45175\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__45178\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10231\ : Odrv4
    port map (
            O => \N__45175\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10230\ : InMux
    port map (
            O => \N__45170\,
            I => \N__45166\
        );

    \I__10229\ : CascadeMux
    port map (
            O => \N__45169\,
            I => \N__45163\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__45166\,
            I => \N__45160\
        );

    \I__10227\ : InMux
    port map (
            O => \N__45163\,
            I => \N__45157\
        );

    \I__10226\ : Span4Mux_h
    port map (
            O => \N__45160\,
            I => \N__45152\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__45157\,
            I => \N__45152\
        );

    \I__10224\ : Span4Mux_v
    port map (
            O => \N__45152\,
            I => \N__45148\
        );

    \I__10223\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45145\
        );

    \I__10222\ : Span4Mux_v
    port map (
            O => \N__45148\,
            I => \N__45141\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__45145\,
            I => \N__45138\
        );

    \I__10220\ : InMux
    port map (
            O => \N__45144\,
            I => \N__45135\
        );

    \I__10219\ : Span4Mux_h
    port map (
            O => \N__45141\,
            I => \N__45132\
        );

    \I__10218\ : Span4Mux_v
    port map (
            O => \N__45138\,
            I => \N__45127\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__45135\,
            I => \N__45127\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__45132\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__45127\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10214\ : InMux
    port map (
            O => \N__45122\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__10213\ : CascadeMux
    port map (
            O => \N__45119\,
            I => \N__45116\
        );

    \I__10212\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45113\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45110\
        );

    \I__10210\ : Odrv4
    port map (
            O => \N__45110\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__10209\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45104\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__45104\,
            I => \N__45101\
        );

    \I__10207\ : Odrv4
    port map (
            O => \N__45101\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__10206\ : CascadeMux
    port map (
            O => \N__45098\,
            I => \N__45084\
        );

    \I__10205\ : CascadeMux
    port map (
            O => \N__45097\,
            I => \N__45080\
        );

    \I__10204\ : CascadeMux
    port map (
            O => \N__45096\,
            I => \N__45076\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__45095\,
            I => \N__45072\
        );

    \I__10202\ : CascadeMux
    port map (
            O => \N__45094\,
            I => \N__45068\
        );

    \I__10201\ : CascadeMux
    port map (
            O => \N__45093\,
            I => \N__45064\
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__45092\,
            I => \N__45060\
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__45091\,
            I => \N__45055\
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__45090\,
            I => \N__45051\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__45089\,
            I => \N__45047\
        );

    \I__10196\ : InMux
    port map (
            O => \N__45088\,
            I => \N__45041\
        );

    \I__10195\ : InMux
    port map (
            O => \N__45087\,
            I => \N__45021\
        );

    \I__10194\ : InMux
    port map (
            O => \N__45084\,
            I => \N__45021\
        );

    \I__10193\ : InMux
    port map (
            O => \N__45083\,
            I => \N__45021\
        );

    \I__10192\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45021\
        );

    \I__10191\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45021\
        );

    \I__10190\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45021\
        );

    \I__10189\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45021\
        );

    \I__10188\ : InMux
    port map (
            O => \N__45072\,
            I => \N__45004\
        );

    \I__10187\ : InMux
    port map (
            O => \N__45071\,
            I => \N__45004\
        );

    \I__10186\ : InMux
    port map (
            O => \N__45068\,
            I => \N__45004\
        );

    \I__10185\ : InMux
    port map (
            O => \N__45067\,
            I => \N__45004\
        );

    \I__10184\ : InMux
    port map (
            O => \N__45064\,
            I => \N__45004\
        );

    \I__10183\ : InMux
    port map (
            O => \N__45063\,
            I => \N__45004\
        );

    \I__10182\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45004\
        );

    \I__10181\ : InMux
    port map (
            O => \N__45059\,
            I => \N__45004\
        );

    \I__10180\ : InMux
    port map (
            O => \N__45058\,
            I => \N__44989\
        );

    \I__10179\ : InMux
    port map (
            O => \N__45055\,
            I => \N__44989\
        );

    \I__10178\ : InMux
    port map (
            O => \N__45054\,
            I => \N__44989\
        );

    \I__10177\ : InMux
    port map (
            O => \N__45051\,
            I => \N__44989\
        );

    \I__10176\ : InMux
    port map (
            O => \N__45050\,
            I => \N__44989\
        );

    \I__10175\ : InMux
    port map (
            O => \N__45047\,
            I => \N__44989\
        );

    \I__10174\ : InMux
    port map (
            O => \N__45046\,
            I => \N__44989\
        );

    \I__10173\ : InMux
    port map (
            O => \N__45045\,
            I => \N__44978\
        );

    \I__10172\ : InMux
    port map (
            O => \N__45044\,
            I => \N__44975\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__45041\,
            I => \N__44972\
        );

    \I__10170\ : InMux
    port map (
            O => \N__45040\,
            I => \N__44969\
        );

    \I__10169\ : CascadeMux
    port map (
            O => \N__45039\,
            I => \N__44966\
        );

    \I__10168\ : CascadeMux
    port map (
            O => \N__45038\,
            I => \N__44962\
        );

    \I__10167\ : CascadeMux
    port map (
            O => \N__45037\,
            I => \N__44958\
        );

    \I__10166\ : CascadeMux
    port map (
            O => \N__45036\,
            I => \N__44954\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__45021\,
            I => \N__44950\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__45004\,
            I => \N__44945\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44989\,
            I => \N__44945\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44988\,
            I => \N__44942\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44987\,
            I => \N__44935\
        );

    \I__10160\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44935\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44985\,
            I => \N__44935\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44926\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44926\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44926\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44981\,
            I => \N__44926\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44978\,
            I => \N__44921\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44975\,
            I => \N__44914\
        );

    \I__10152\ : Span4Mux_s1_v
    port map (
            O => \N__44972\,
            I => \N__44914\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__44969\,
            I => \N__44914\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44966\,
            I => \N__44897\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44897\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44962\,
            I => \N__44897\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44897\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44897\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44897\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44897\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44897\
        );

    \I__10142\ : Span4Mux_v
    port map (
            O => \N__44950\,
            I => \N__44892\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__44945\,
            I => \N__44892\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44942\,
            I => \N__44883\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44935\,
            I => \N__44883\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44926\,
            I => \N__44883\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44880\
        );

    \I__10136\ : CascadeMux
    port map (
            O => \N__44924\,
            I => \N__44869\
        );

    \I__10135\ : Span12Mux_s5_v
    port map (
            O => \N__44921\,
            I => \N__44865\
        );

    \I__10134\ : Span4Mux_h
    port map (
            O => \N__44914\,
            I => \N__44862\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44897\,
            I => \N__44859\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__44892\,
            I => \N__44856\
        );

    \I__10131\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44851\
        );

    \I__10130\ : InMux
    port map (
            O => \N__44890\,
            I => \N__44851\
        );

    \I__10129\ : Span4Mux_v
    port map (
            O => \N__44883\,
            I => \N__44848\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__44880\,
            I => \N__44845\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44838\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44838\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44838\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44876\,
            I => \N__44829\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44875\,
            I => \N__44829\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44829\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44873\,
            I => \N__44829\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44822\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44822\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44868\,
            I => \N__44822\
        );

    \I__10117\ : Span12Mux_v
    port map (
            O => \N__44865\,
            I => \N__44819\
        );

    \I__10116\ : Sp12to4
    port map (
            O => \N__44862\,
            I => \N__44816\
        );

    \I__10115\ : Span12Mux_s9_h
    port map (
            O => \N__44859\,
            I => \N__44809\
        );

    \I__10114\ : Sp12to4
    port map (
            O => \N__44856\,
            I => \N__44809\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44851\,
            I => \N__44809\
        );

    \I__10112\ : Span4Mux_v
    port map (
            O => \N__44848\,
            I => \N__44800\
        );

    \I__10111\ : Span4Mux_v
    port map (
            O => \N__44845\,
            I => \N__44800\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__44838\,
            I => \N__44800\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44829\,
            I => \N__44800\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__44822\,
            I => \N__44797\
        );

    \I__10107\ : Span12Mux_h
    port map (
            O => \N__44819\,
            I => \N__44794\
        );

    \I__10106\ : Span12Mux_s10_v
    port map (
            O => \N__44816\,
            I => \N__44789\
        );

    \I__10105\ : Span12Mux_h
    port map (
            O => \N__44809\,
            I => \N__44789\
        );

    \I__10104\ : Span4Mux_h
    port map (
            O => \N__44800\,
            I => \N__44786\
        );

    \I__10103\ : Span4Mux_v
    port map (
            O => \N__44797\,
            I => \N__44783\
        );

    \I__10102\ : Odrv12
    port map (
            O => \N__44794\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10101\ : Odrv12
    port map (
            O => \N__44789\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__44786\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10099\ : Odrv4
    port map (
            O => \N__44783\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10098\ : CascadeMux
    port map (
            O => \N__44774\,
            I => \N__44771\
        );

    \I__10097\ : InMux
    port map (
            O => \N__44771\,
            I => \N__44768\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44768\,
            I => \N__44765\
        );

    \I__10095\ : Span4Mux_v
    port map (
            O => \N__44765\,
            I => \N__44762\
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__44762\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44747\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44758\,
            I => \N__44747\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44736\
        );

    \I__10090\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44736\
        );

    \I__10089\ : InMux
    port map (
            O => \N__44755\,
            I => \N__44736\
        );

    \I__10088\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44736\
        );

    \I__10087\ : InMux
    port map (
            O => \N__44753\,
            I => \N__44736\
        );

    \I__10086\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44701\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__44747\,
            I => \N__44696\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44736\,
            I => \N__44696\
        );

    \I__10083\ : InMux
    port map (
            O => \N__44735\,
            I => \N__44679\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44679\
        );

    \I__10081\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44679\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44679\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44731\,
            I => \N__44679\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44730\,
            I => \N__44679\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44729\,
            I => \N__44679\
        );

    \I__10076\ : InMux
    port map (
            O => \N__44728\,
            I => \N__44679\
        );

    \I__10075\ : InMux
    port map (
            O => \N__44727\,
            I => \N__44674\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44726\,
            I => \N__44669\
        );

    \I__10073\ : InMux
    port map (
            O => \N__44725\,
            I => \N__44669\
        );

    \I__10072\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44642\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44723\,
            I => \N__44642\
        );

    \I__10070\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44642\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44642\
        );

    \I__10068\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44642\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44642\
        );

    \I__10066\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44642\
        );

    \I__10065\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44625\
        );

    \I__10064\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44625\
        );

    \I__10063\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44625\
        );

    \I__10062\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44625\
        );

    \I__10061\ : InMux
    port map (
            O => \N__44713\,
            I => \N__44625\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44712\,
            I => \N__44625\
        );

    \I__10059\ : InMux
    port map (
            O => \N__44711\,
            I => \N__44625\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44710\,
            I => \N__44625\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44709\,
            I => \N__44609\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44609\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44609\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44609\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44705\,
            I => \N__44609\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44606\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44701\,
            I => \N__44599\
        );

    \I__10050\ : Span4Mux_h
    port map (
            O => \N__44696\,
            I => \N__44599\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__44679\,
            I => \N__44599\
        );

    \I__10048\ : InMux
    port map (
            O => \N__44678\,
            I => \N__44586\
        );

    \I__10047\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44586\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__44674\,
            I => \N__44581\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__44669\,
            I => \N__44581\
        );

    \I__10044\ : InMux
    port map (
            O => \N__44668\,
            I => \N__44564\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44564\
        );

    \I__10042\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44564\
        );

    \I__10041\ : InMux
    port map (
            O => \N__44665\,
            I => \N__44564\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44664\,
            I => \N__44564\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44564\
        );

    \I__10038\ : InMux
    port map (
            O => \N__44662\,
            I => \N__44564\
        );

    \I__10037\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44564\
        );

    \I__10036\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44557\
        );

    \I__10035\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44557\
        );

    \I__10034\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44557\
        );

    \I__10033\ : CascadeMux
    port map (
            O => \N__44657\,
            I => \N__44553\
        );

    \I__10032\ : LocalMux
    port map (
            O => \N__44642\,
            I => \N__44545\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__44625\,
            I => \N__44545\
        );

    \I__10030\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44534\
        );

    \I__10029\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44534\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44534\
        );

    \I__10027\ : InMux
    port map (
            O => \N__44621\,
            I => \N__44534\
        );

    \I__10026\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44534\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__44609\,
            I => \N__44527\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__44606\,
            I => \N__44527\
        );

    \I__10023\ : Span4Mux_v
    port map (
            O => \N__44599\,
            I => \N__44527\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44598\,
            I => \N__44510\
        );

    \I__10021\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44510\
        );

    \I__10020\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44510\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44595\,
            I => \N__44510\
        );

    \I__10018\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44510\
        );

    \I__10017\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44510\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44592\,
            I => \N__44510\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44591\,
            I => \N__44510\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__44586\,
            I => \N__44507\
        );

    \I__10013\ : Span4Mux_h
    port map (
            O => \N__44581\,
            I => \N__44500\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44500\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44557\,
            I => \N__44500\
        );

    \I__10010\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44489\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44489\
        );

    \I__10008\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44489\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44489\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44550\,
            I => \N__44489\
        );

    \I__10005\ : Odrv12
    port map (
            O => \N__44545\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44534\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10003\ : Odrv4
    port map (
            O => \N__44527\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__44510\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10001\ : Odrv4
    port map (
            O => \N__44507\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10000\ : Odrv4
    port map (
            O => \N__44500\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__44489\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__9998\ : InMux
    port map (
            O => \N__44474\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44471\,
            I => \N__44456\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44470\,
            I => \N__44456\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44439\
        );

    \I__9994\ : InMux
    port map (
            O => \N__44468\,
            I => \N__44439\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44467\,
            I => \N__44439\
        );

    \I__9992\ : InMux
    port map (
            O => \N__44466\,
            I => \N__44439\
        );

    \I__9991\ : InMux
    port map (
            O => \N__44465\,
            I => \N__44439\
        );

    \I__9990\ : InMux
    port map (
            O => \N__44464\,
            I => \N__44439\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44463\,
            I => \N__44439\
        );

    \I__9988\ : InMux
    port map (
            O => \N__44462\,
            I => \N__44439\
        );

    \I__9987\ : InMux
    port map (
            O => \N__44461\,
            I => \N__44436\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__44456\,
            I => \N__44433\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__44439\,
            I => \N__44430\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44436\,
            I => \N__44421\
        );

    \I__9983\ : Span4Mux_h
    port map (
            O => \N__44433\,
            I => \N__44421\
        );

    \I__9982\ : Span4Mux_h
    port map (
            O => \N__44430\,
            I => \N__44418\
        );

    \I__9981\ : InMux
    port map (
            O => \N__44429\,
            I => \N__44409\
        );

    \I__9980\ : InMux
    port map (
            O => \N__44428\,
            I => \N__44409\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44409\
        );

    \I__9978\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44409\
        );

    \I__9977\ : Span4Mux_h
    port map (
            O => \N__44421\,
            I => \N__44406\
        );

    \I__9976\ : Span4Mux_h
    port map (
            O => \N__44418\,
            I => \N__44403\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__44409\,
            I => \N__44400\
        );

    \I__9974\ : Odrv4
    port map (
            O => \N__44406\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9973\ : Odrv4
    port map (
            O => \N__44403\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9972\ : Odrv12
    port map (
            O => \N__44400\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44389\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44386\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__44389\,
            I => \N__44382\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__44386\,
            I => \N__44379\
        );

    \I__9967\ : InMux
    port map (
            O => \N__44385\,
            I => \N__44376\
        );

    \I__9966\ : Span4Mux_v
    port map (
            O => \N__44382\,
            I => \N__44371\
        );

    \I__9965\ : Span4Mux_h
    port map (
            O => \N__44379\,
            I => \N__44371\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__44376\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9963\ : Odrv4
    port map (
            O => \N__44371\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9962\ : CascadeMux
    port map (
            O => \N__44366\,
            I => \N__44363\
        );

    \I__9961\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44357\
        );

    \I__9960\ : InMux
    port map (
            O => \N__44362\,
            I => \N__44357\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__44357\,
            I => \N__44352\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44349\
        );

    \I__9957\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44346\
        );

    \I__9956\ : Span4Mux_h
    port map (
            O => \N__44352\,
            I => \N__44339\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__44349\,
            I => \N__44339\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44339\
        );

    \I__9953\ : Odrv4
    port map (
            O => \N__44339\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44332\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44329\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__44332\,
            I => \N__44325\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__44329\,
            I => \N__44322\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44319\
        );

    \I__9947\ : Span4Mux_h
    port map (
            O => \N__44325\,
            I => \N__44316\
        );

    \I__9946\ : Odrv12
    port map (
            O => \N__44322\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__44319\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9944\ : Odrv4
    port map (
            O => \N__44316\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__44309\,
            I => \N__44306\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44306\,
            I => \N__44302\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44305\,
            I => \N__44299\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44302\,
            I => \N__44295\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44292\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44289\
        );

    \I__9937\ : Span4Mux_v
    port map (
            O => \N__44295\,
            I => \N__44285\
        );

    \I__9936\ : Span4Mux_v
    port map (
            O => \N__44292\,
            I => \N__44280\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__44289\,
            I => \N__44280\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44288\,
            I => \N__44277\
        );

    \I__9933\ : Span4Mux_h
    port map (
            O => \N__44285\,
            I => \N__44274\
        );

    \I__9932\ : Span4Mux_h
    port map (
            O => \N__44280\,
            I => \N__44269\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__44277\,
            I => \N__44269\
        );

    \I__9930\ : Odrv4
    port map (
            O => \N__44274\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__44269\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9928\ : InMux
    port map (
            O => \N__44264\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__9927\ : CascadeMux
    port map (
            O => \N__44261\,
            I => \N__44257\
        );

    \I__9926\ : CascadeMux
    port map (
            O => \N__44260\,
            I => \N__44254\
        );

    \I__9925\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44249\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44254\,
            I => \N__44249\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__44249\,
            I => \N__44245\
        );

    \I__9922\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44242\
        );

    \I__9921\ : Span12Mux_s10_h
    port map (
            O => \N__44245\,
            I => \N__44239\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__44242\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9919\ : Odrv12
    port map (
            O => \N__44239\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9918\ : CascadeMux
    port map (
            O => \N__44234\,
            I => \N__44231\
        );

    \I__9917\ : InMux
    port map (
            O => \N__44231\,
            I => \N__44227\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44230\,
            I => \N__44224\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__44227\,
            I => \N__44219\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__44224\,
            I => \N__44216\
        );

    \I__9913\ : CascadeMux
    port map (
            O => \N__44223\,
            I => \N__44213\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44222\,
            I => \N__44210\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__44219\,
            I => \N__44205\
        );

    \I__9910\ : Span4Mux_v
    port map (
            O => \N__44216\,
            I => \N__44205\
        );

    \I__9909\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44202\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__44210\,
            I => \N__44199\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__44205\,
            I => \N__44196\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__44202\,
            I => \N__44191\
        );

    \I__9905\ : Span4Mux_h
    port map (
            O => \N__44199\,
            I => \N__44191\
        );

    \I__9904\ : Odrv4
    port map (
            O => \N__44196\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__44191\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9902\ : InMux
    port map (
            O => \N__44186\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__9901\ : CascadeMux
    port map (
            O => \N__44183\,
            I => \N__44179\
        );

    \I__9900\ : CascadeMux
    port map (
            O => \N__44182\,
            I => \N__44176\
        );

    \I__9899\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44171\
        );

    \I__9898\ : InMux
    port map (
            O => \N__44176\,
            I => \N__44171\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__44171\,
            I => \N__44167\
        );

    \I__9896\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44164\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__44167\,
            I => \N__44161\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__44164\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9893\ : Odrv4
    port map (
            O => \N__44161\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9892\ : CascadeMux
    port map (
            O => \N__44156\,
            I => \N__44152\
        );

    \I__9891\ : CascadeMux
    port map (
            O => \N__44155\,
            I => \N__44149\
        );

    \I__9890\ : InMux
    port map (
            O => \N__44152\,
            I => \N__44146\
        );

    \I__9889\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44143\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__44146\,
            I => \N__44138\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__44143\,
            I => \N__44138\
        );

    \I__9886\ : Span4Mux_h
    port map (
            O => \N__44138\,
            I => \N__44133\
        );

    \I__9885\ : InMux
    port map (
            O => \N__44137\,
            I => \N__44130\
        );

    \I__9884\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44127\
        );

    \I__9883\ : Span4Mux_v
    port map (
            O => \N__44133\,
            I => \N__44124\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__44130\,
            I => \N__44119\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__44127\,
            I => \N__44119\
        );

    \I__9880\ : Odrv4
    port map (
            O => \N__44124\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__44119\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9878\ : InMux
    port map (
            O => \N__44114\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__9877\ : CascadeMux
    port map (
            O => \N__44111\,
            I => \N__44108\
        );

    \I__9876\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44105\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__44105\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__9874\ : InMux
    port map (
            O => \N__44102\,
            I => \N__44099\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__44099\,
            I => \N__44096\
        );

    \I__9872\ : Odrv4
    port map (
            O => \N__44096\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__9871\ : CascadeMux
    port map (
            O => \N__44093\,
            I => \N__44090\
        );

    \I__9870\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44087\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__44087\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__9868\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44081\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__44081\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__9866\ : CascadeMux
    port map (
            O => \N__44078\,
            I => \N__44075\
        );

    \I__9865\ : InMux
    port map (
            O => \N__44075\,
            I => \N__44072\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__44072\,
            I => \N__44069\
        );

    \I__9863\ : Span12Mux_s9_h
    port map (
            O => \N__44069\,
            I => \N__44066\
        );

    \I__9862\ : Odrv12
    port map (
            O => \N__44066\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__9861\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44060\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__44060\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__9859\ : CascadeMux
    port map (
            O => \N__44057\,
            I => \N__44054\
        );

    \I__9858\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44051\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__44051\,
            I => \N__44048\
        );

    \I__9856\ : Span4Mux_h
    port map (
            O => \N__44048\,
            I => \N__44045\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__44045\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__9854\ : InMux
    port map (
            O => \N__44042\,
            I => \N__44039\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__44039\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__44036\,
            I => \N__44033\
        );

    \I__9851\ : InMux
    port map (
            O => \N__44033\,
            I => \N__44030\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__44030\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__9849\ : InMux
    port map (
            O => \N__44027\,
            I => \N__44024\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__44024\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__9847\ : CascadeMux
    port map (
            O => \N__44021\,
            I => \N__44018\
        );

    \I__9846\ : InMux
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__44015\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__9844\ : InMux
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__44009\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__9842\ : CascadeMux
    port map (
            O => \N__44006\,
            I => \N__44003\
        );

    \I__9841\ : InMux
    port map (
            O => \N__44003\,
            I => \N__44000\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__44000\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43994\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43994\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__9837\ : CascadeMux
    port map (
            O => \N__43991\,
            I => \N__43988\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43988\,
            I => \N__43985\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43985\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43982\,
            I => \N__43979\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43979\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__43976\,
            I => \N__43973\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43970\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__43970\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43964\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43964\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__9827\ : CascadeMux
    port map (
            O => \N__43961\,
            I => \N__43958\
        );

    \I__9826\ : InMux
    port map (
            O => \N__43958\,
            I => \N__43955\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__43955\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43949\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43949\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__43946\,
            I => \N__43943\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43943\,
            I => \N__43940\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__43940\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__43937\,
            I => \N__43934\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43934\,
            I => \N__43931\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43931\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43928\,
            I => \N__43925\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43925\,
            I => \N__43922\
        );

    \I__9814\ : Span4Mux_h
    port map (
            O => \N__43922\,
            I => \N__43919\
        );

    \I__9813\ : Span4Mux_h
    port map (
            O => \N__43919\,
            I => \N__43916\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__43916\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__9811\ : CascadeMux
    port map (
            O => \N__43913\,
            I => \N__43910\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43910\,
            I => \N__43907\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43907\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43904\,
            I => \N__43901\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43901\,
            I => \N__43898\
        );

    \I__9806\ : Odrv12
    port map (
            O => \N__43898\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__9805\ : InMux
    port map (
            O => \N__43895\,
            I => \N__43889\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43894\,
            I => \N__43884\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43893\,
            I => \N__43884\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43892\,
            I => \N__43881\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__43889\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__43884\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43881\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9798\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43870\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43873\,
            I => \N__43867\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43863\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__43867\,
            I => \N__43859\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43866\,
            I => \N__43856\
        );

    \I__9793\ : Span4Mux_h
    port map (
            O => \N__43863\,
            I => \N__43853\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43850\
        );

    \I__9791\ : Odrv12
    port map (
            O => \N__43859\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__43856\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__43853\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__43850\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9787\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43837\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43833\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__43837\,
            I => \N__43830\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43827\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43833\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__9782\ : Odrv12
    port map (
            O => \N__43830\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43827\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43817\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43817\,
            I => \N__43814\
        );

    \I__9778\ : Span12Mux_v
    port map (
            O => \N__43814\,
            I => \N__43811\
        );

    \I__9777\ : Odrv12
    port map (
            O => \N__43811\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__9776\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43804\
        );

    \I__9775\ : InMux
    port map (
            O => \N__43807\,
            I => \N__43801\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43795\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43801\,
            I => \N__43792\
        );

    \I__9772\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43789\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43784\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43798\,
            I => \N__43784\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__43795\,
            I => \N__43781\
        );

    \I__9768\ : Odrv12
    port map (
            O => \N__43792\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43789\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__43784\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__9765\ : Odrv4
    port map (
            O => \N__43781\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__9764\ : CascadeMux
    port map (
            O => \N__43772\,
            I => \N__43769\
        );

    \I__9763\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43766\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43766\,
            I => \N__43762\
        );

    \I__9761\ : InMux
    port map (
            O => \N__43765\,
            I => \N__43759\
        );

    \I__9760\ : Span4Mux_h
    port map (
            O => \N__43762\,
            I => \N__43756\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43759\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__43756\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__9757\ : CascadeMux
    port map (
            O => \N__43751\,
            I => \N__43748\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43748\,
            I => \N__43745\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__43745\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43742\,
            I => \N__43739\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43739\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__9752\ : CascadeMux
    port map (
            O => \N__43736\,
            I => \N__43731\
        );

    \I__9751\ : CascadeMux
    port map (
            O => \N__43735\,
            I => \N__43728\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43734\,
            I => \N__43720\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43731\,
            I => \N__43720\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43720\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43727\,
            I => \N__43717\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__43720\,
            I => \N__43714\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__43717\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__9744\ : Odrv4
    port map (
            O => \N__43714\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43709\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43706\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__9741\ : CascadeMux
    port map (
            O => \N__43703\,
            I => \N__43700\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43691\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43699\,
            I => \N__43691\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43698\,
            I => \N__43691\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43691\,
            I => \N__43687\
        );

    \I__9736\ : InMux
    port map (
            O => \N__43690\,
            I => \N__43684\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__43687\,
            I => \N__43681\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43684\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__43681\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__9732\ : CascadeMux
    port map (
            O => \N__43676\,
            I => \N__43673\
        );

    \I__9731\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43670\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__43670\,
            I => \N__43667\
        );

    \I__9729\ : Span4Mux_v
    port map (
            O => \N__43667\,
            I => \N__43664\
        );

    \I__9728\ : Odrv4
    port map (
            O => \N__43664\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__9727\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43656\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43651\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43659\,
            I => \N__43651\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__43656\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__43651\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__9722\ : CascadeMux
    port map (
            O => \N__43646\,
            I => \N__43643\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43643\,
            I => \N__43636\
        );

    \I__9720\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43636\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43633\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__43636\,
            I => \N__43630\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43633\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__9716\ : Odrv4
    port map (
            O => \N__43630\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__9715\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43622\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__43622\,
            I => \N__43619\
        );

    \I__9713\ : Odrv12
    port map (
            O => \N__43619\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__9712\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43609\
        );

    \I__9710\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43606\
        );

    \I__9709\ : Odrv4
    port map (
            O => \N__43609\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43606\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__9707\ : CascadeMux
    port map (
            O => \N__43601\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\
        );

    \I__9706\ : CascadeMux
    port map (
            O => \N__43598\,
            I => \N__43595\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43595\,
            I => \N__43589\
        );

    \I__9704\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43589\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__43589\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__9702\ : InMux
    port map (
            O => \N__43586\,
            I => \N__43580\
        );

    \I__9701\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43577\
        );

    \I__9700\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43574\
        );

    \I__9699\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43571\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__43580\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__43577\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__43574\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__43571\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9694\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43559\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__43559\,
            I => \N__43555\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43551\
        );

    \I__9691\ : Span4Mux_h
    port map (
            O => \N__43555\,
            I => \N__43548\
        );

    \I__9690\ : InMux
    port map (
            O => \N__43554\,
            I => \N__43545\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__43551\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__9688\ : Odrv4
    port map (
            O => \N__43548\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__43545\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__9686\ : InMux
    port map (
            O => \N__43538\,
            I => \N__43532\
        );

    \I__9685\ : InMux
    port map (
            O => \N__43537\,
            I => \N__43532\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__43532\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43526\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43526\,
            I => \N__43521\
        );

    \I__9681\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43516\
        );

    \I__9680\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43516\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__43521\,
            I => \N__43512\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43516\,
            I => \N__43509\
        );

    \I__9677\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43506\
        );

    \I__9676\ : Odrv4
    port map (
            O => \N__43512\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9675\ : Odrv12
    port map (
            O => \N__43509\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__43506\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43494\
        );

    \I__9672\ : InMux
    port map (
            O => \N__43498\,
            I => \N__43489\
        );

    \I__9671\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43489\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43494\,
            I => \N__43486\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__43489\,
            I => \N__43483\
        );

    \I__9668\ : Span4Mux_v
    port map (
            O => \N__43486\,
            I => \N__43479\
        );

    \I__9667\ : Span4Mux_v
    port map (
            O => \N__43483\,
            I => \N__43476\
        );

    \I__9666\ : InMux
    port map (
            O => \N__43482\,
            I => \N__43473\
        );

    \I__9665\ : Odrv4
    port map (
            O => \N__43479\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9664\ : Odrv4
    port map (
            O => \N__43476\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__43473\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9662\ : InMux
    port map (
            O => \N__43466\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__9661\ : CascadeMux
    port map (
            O => \N__43463\,
            I => \N__43458\
        );

    \I__9660\ : InMux
    port map (
            O => \N__43462\,
            I => \N__43455\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43461\,
            I => \N__43450\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43458\,
            I => \N__43450\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__43455\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__43450\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43445\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__9654\ : CascadeMux
    port map (
            O => \N__43442\,
            I => \N__43437\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43434\
        );

    \I__9652\ : InMux
    port map (
            O => \N__43440\,
            I => \N__43429\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43437\,
            I => \N__43429\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__43434\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__43429\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__9648\ : InMux
    port map (
            O => \N__43424\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__9647\ : InMux
    port map (
            O => \N__43421\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43418\,
            I => \bfn_17_21_0_\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43415\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__9644\ : InMux
    port map (
            O => \N__43412\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__9643\ : InMux
    port map (
            O => \N__43409\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43406\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43399\
        );

    \I__9640\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43396\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__43399\,
            I => \N__43393\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__43396\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__9637\ : Odrv4
    port map (
            O => \N__43393\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43388\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__9635\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43381\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43384\,
            I => \N__43378\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43375\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__43378\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__9631\ : Odrv4
    port map (
            O => \N__43375\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43370\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43363\
        );

    \I__9628\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43360\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43363\,
            I => \N__43357\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__43360\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__9625\ : Odrv4
    port map (
            O => \N__43357\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__9624\ : InMux
    port map (
            O => \N__43352\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43349\,
            I => \N__43346\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__43346\,
            I => \N__43342\
        );

    \I__9621\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43339\
        );

    \I__9620\ : Span4Mux_v
    port map (
            O => \N__43342\,
            I => \N__43336\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__43339\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__43336\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43331\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43328\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__9615\ : InMux
    port map (
            O => \N__43325\,
            I => \bfn_17_20_0_\
        );

    \I__9614\ : InMux
    port map (
            O => \N__43322\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__9613\ : InMux
    port map (
            O => \N__43319\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__9612\ : InMux
    port map (
            O => \N__43316\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__9611\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43309\
        );

    \I__9610\ : InMux
    port map (
            O => \N__43312\,
            I => \N__43306\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__43309\,
            I => \N__43303\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__43306\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__43303\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__9606\ : InMux
    port map (
            O => \N__43298\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__9605\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43291\
        );

    \I__9604\ : InMux
    port map (
            O => \N__43294\,
            I => \N__43288\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__43291\,
            I => \N__43285\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__43288\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__9601\ : Odrv4
    port map (
            O => \N__43285\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__9600\ : InMux
    port map (
            O => \N__43280\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__9599\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43273\
        );

    \I__9598\ : InMux
    port map (
            O => \N__43276\,
            I => \N__43270\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__43273\,
            I => \N__43267\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__43270\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__9595\ : Odrv4
    port map (
            O => \N__43267\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__9594\ : InMux
    port map (
            O => \N__43262\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43259\,
            I => \N__43255\
        );

    \I__9592\ : InMux
    port map (
            O => \N__43258\,
            I => \N__43252\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__43255\,
            I => \N__43249\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43252\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__9589\ : Odrv12
    port map (
            O => \N__43249\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43244\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__9587\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43237\
        );

    \I__9586\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43234\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43237\,
            I => \N__43231\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__43234\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__9583\ : Odrv12
    port map (
            O => \N__43231\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__9582\ : InMux
    port map (
            O => \N__43226\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__9581\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43219\
        );

    \I__9580\ : InMux
    port map (
            O => \N__43222\,
            I => \N__43216\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__43219\,
            I => \N__43213\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__43216\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__9577\ : Odrv4
    port map (
            O => \N__43213\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__9576\ : InMux
    port map (
            O => \N__43208\,
            I => \bfn_17_19_0_\
        );

    \I__9575\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43202\,
            I => \N__43198\
        );

    \I__9573\ : InMux
    port map (
            O => \N__43201\,
            I => \N__43195\
        );

    \I__9572\ : Span4Mux_h
    port map (
            O => \N__43198\,
            I => \N__43192\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__43195\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__43192\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__9569\ : InMux
    port map (
            O => \N__43187\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__9568\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43180\
        );

    \I__9567\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43177\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43174\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__43177\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__9564\ : Odrv4
    port map (
            O => \N__43174\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__9563\ : InMux
    port map (
            O => \N__43169\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__9562\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43163\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43163\,
            I => \N__43160\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__43160\,
            I => \N__43157\
        );

    \I__9559\ : Odrv4
    port map (
            O => \N__43157\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__9558\ : CascadeMux
    port map (
            O => \N__43154\,
            I => \N__43151\
        );

    \I__9557\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43148\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__43148\,
            I => \N__43145\
        );

    \I__9555\ : Span4Mux_v
    port map (
            O => \N__43145\,
            I => \N__43142\
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__43142\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__9553\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43136\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__43136\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__9551\ : CascadeMux
    port map (
            O => \N__43133\,
            I => \N__43130\
        );

    \I__9550\ : InMux
    port map (
            O => \N__43130\,
            I => \N__43127\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__43127\,
            I => \N__43123\
        );

    \I__9548\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43120\
        );

    \I__9547\ : Odrv4
    port map (
            O => \N__43123\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__43120\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__9545\ : InMux
    port map (
            O => \N__43115\,
            I => \N__43112\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__43112\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__9543\ : InMux
    port map (
            O => \N__43109\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28\
        );

    \I__9542\ : InMux
    port map (
            O => \N__43106\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__9541\ : InMux
    port map (
            O => \N__43103\,
            I => \N__43099\
        );

    \I__9540\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43096\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__43099\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__43096\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__9537\ : CascadeMux
    port map (
            O => \N__43091\,
            I => \N__43087\
        );

    \I__9536\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43084\
        );

    \I__9535\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43080\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__43084\,
            I => \N__43077\
        );

    \I__9533\ : InMux
    port map (
            O => \N__43083\,
            I => \N__43074\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__43080\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9531\ : Odrv4
    port map (
            O => \N__43077\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__43074\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9529\ : CascadeMux
    port map (
            O => \N__43067\,
            I => \N__43064\
        );

    \I__9528\ : InMux
    port map (
            O => \N__43064\,
            I => \N__43061\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__43061\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__9526\ : InMux
    port map (
            O => \N__43058\,
            I => \N__43054\
        );

    \I__9525\ : InMux
    port map (
            O => \N__43057\,
            I => \N__43051\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__43054\,
            I => \N__43048\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__43051\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__9522\ : Odrv4
    port map (
            O => \N__43048\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__9521\ : InMux
    port map (
            O => \N__43043\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__9520\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__43037\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__43034\,
            I => \N__43030\
        );

    \I__9517\ : InMux
    port map (
            O => \N__43033\,
            I => \N__43027\
        );

    \I__9516\ : InMux
    port map (
            O => \N__43030\,
            I => \N__43024\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__43027\,
            I => \N__43021\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__43024\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__43021\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__9512\ : InMux
    port map (
            O => \N__43016\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__9511\ : InMux
    port map (
            O => \N__43013\,
            I => \N__43010\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__43007\,
            I => \N__43004\
        );

    \I__9508\ : Odrv4
    port map (
            O => \N__43004\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__9507\ : CascadeMux
    port map (
            O => \N__43001\,
            I => \N__42998\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42998\,
            I => \N__42995\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__42995\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42992\,
            I => \N__42989\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__42989\,
            I => \N__42986\
        );

    \I__9502\ : Span4Mux_v
    port map (
            O => \N__42986\,
            I => \N__42983\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__42983\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__9500\ : CascadeMux
    port map (
            O => \N__42980\,
            I => \N__42977\
        );

    \I__9499\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42974\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42974\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__42971\,
            I => \N__42968\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42965\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42965\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__9494\ : CascadeMux
    port map (
            O => \N__42962\,
            I => \N__42959\
        );

    \I__9493\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42956\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__42956\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42950\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__42950\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42944\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__42944\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__9487\ : CascadeMux
    port map (
            O => \N__42941\,
            I => \N__42938\
        );

    \I__9486\ : InMux
    port map (
            O => \N__42938\,
            I => \N__42935\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__42935\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42932\,
            I => \N__42929\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42929\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__9482\ : CascadeMux
    port map (
            O => \N__42926\,
            I => \N__42923\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42923\,
            I => \N__42920\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42920\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42917\,
            I => \N__42914\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__42914\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__9477\ : CascadeMux
    port map (
            O => \N__42911\,
            I => \N__42908\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42905\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42902\,
            I => \N__42899\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__42899\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__9472\ : CascadeMux
    port map (
            O => \N__42896\,
            I => \N__42893\
        );

    \I__9471\ : InMux
    port map (
            O => \N__42893\,
            I => \N__42890\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__42890\,
            I => \N__42887\
        );

    \I__9469\ : Odrv4
    port map (
            O => \N__42887\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__9468\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42881\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42878\
        );

    \I__9466\ : Span4Mux_h
    port map (
            O => \N__42878\,
            I => \N__42875\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__42875\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42866\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42866\,
            I => \N__42863\
        );

    \I__9461\ : Odrv4
    port map (
            O => \N__42863\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__9460\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42857\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42857\,
            I => \N__42854\
        );

    \I__9458\ : Span4Mux_h
    port map (
            O => \N__42854\,
            I => \N__42851\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__42851\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__42848\,
            I => \N__42845\
        );

    \I__9455\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42842\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__42842\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42836\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42836\,
            I => \N__42833\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__42833\,
            I => \N__42830\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__42830\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__9449\ : CascadeMux
    port map (
            O => \N__42827\,
            I => \N__42824\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42821\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42821\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42815\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42815\,
            I => \N__42812\
        );

    \I__9444\ : Odrv4
    port map (
            O => \N__42812\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42806\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__42806\,
            I => \N__42803\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__42803\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42797\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__42797\,
            I => \N__42794\
        );

    \I__9438\ : Odrv4
    port map (
            O => \N__42794\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9437\ : CascadeMux
    port map (
            O => \N__42791\,
            I => \N__42788\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42785\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42785\,
            I => \N__42782\
        );

    \I__9434\ : Odrv4
    port map (
            O => \N__42782\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__9433\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42776\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__42776\,
            I => \N__42773\
        );

    \I__9431\ : Span4Mux_h
    port map (
            O => \N__42773\,
            I => \N__42770\
        );

    \I__9430\ : Odrv4
    port map (
            O => \N__42770\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42767\,
            I => \N__42764\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__42764\,
            I => \N__42761\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__42761\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42758\,
            I => \N__42754\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42757\,
            I => \N__42750\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__42754\,
            I => \N__42746\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42743\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__42750\,
            I => \N__42740\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42737\
        );

    \I__9420\ : Span4Mux_v
    port map (
            O => \N__42746\,
            I => \N__42734\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__42743\,
            I => \N__42731\
        );

    \I__9418\ : Span4Mux_v
    port map (
            O => \N__42740\,
            I => \N__42726\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__42737\,
            I => \N__42726\
        );

    \I__9416\ : Span4Mux_h
    port map (
            O => \N__42734\,
            I => \N__42723\
        );

    \I__9415\ : Span4Mux_v
    port map (
            O => \N__42731\,
            I => \N__42720\
        );

    \I__9414\ : Span4Mux_h
    port map (
            O => \N__42726\,
            I => \N__42715\
        );

    \I__9413\ : Span4Mux_h
    port map (
            O => \N__42723\,
            I => \N__42715\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__42720\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9411\ : Odrv4
    port map (
            O => \N__42715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9410\ : CascadeMux
    port map (
            O => \N__42710\,
            I => \N__42707\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42704\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42701\
        );

    \I__9407\ : Span4Mux_v
    port map (
            O => \N__42701\,
            I => \N__42698\
        );

    \I__9406\ : Span4Mux_h
    port map (
            O => \N__42698\,
            I => \N__42695\
        );

    \I__9405\ : Span4Mux_h
    port map (
            O => \N__42695\,
            I => \N__42692\
        );

    \I__9404\ : Odrv4
    port map (
            O => \N__42692\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__9403\ : CascadeMux
    port map (
            O => \N__42689\,
            I => \N__42686\
        );

    \I__9402\ : InMux
    port map (
            O => \N__42686\,
            I => \N__42683\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__42683\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__9400\ : CascadeMux
    port map (
            O => \N__42680\,
            I => \N__42677\
        );

    \I__9399\ : InMux
    port map (
            O => \N__42677\,
            I => \N__42674\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__42674\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42668\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__42668\,
            I => \N__42665\
        );

    \I__9395\ : Odrv4
    port map (
            O => \N__42665\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9394\ : CascadeMux
    port map (
            O => \N__42662\,
            I => \N__42659\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42659\,
            I => \N__42656\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__42656\,
            I => \N__42653\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__42653\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__9390\ : InMux
    port map (
            O => \N__42650\,
            I => \N__42647\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__9388\ : Odrv4
    port map (
            O => \N__42644\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__42638\,
            I => \N__42635\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__42635\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__9384\ : CascadeMux
    port map (
            O => \N__42632\,
            I => \N__42629\
        );

    \I__9383\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42626\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__42626\,
            I => \N__42623\
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__42623\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42617\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42617\,
            I => \N__42614\
        );

    \I__9378\ : Span4Mux_v
    port map (
            O => \N__42614\,
            I => \N__42611\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__42611\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9376\ : CascadeMux
    port map (
            O => \N__42608\,
            I => \N__42605\
        );

    \I__9375\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42602\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__42602\,
            I => \N__42599\
        );

    \I__9373\ : Odrv4
    port map (
            O => \N__42599\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__9372\ : InMux
    port map (
            O => \N__42596\,
            I => \N__42593\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42593\,
            I => \N__42590\
        );

    \I__9370\ : Span4Mux_h
    port map (
            O => \N__42590\,
            I => \N__42587\
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__42587\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42584\,
            I => \N__42581\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42581\,
            I => \N__42578\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__42578\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9365\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42572\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__42572\,
            I => \N__42567\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42564\
        );

    \I__9362\ : InMux
    port map (
            O => \N__42570\,
            I => \N__42561\
        );

    \I__9361\ : Span4Mux_v
    port map (
            O => \N__42567\,
            I => \N__42556\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__42564\,
            I => \N__42556\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__42561\,
            I => \N__42553\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__42556\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9357\ : Odrv4
    port map (
            O => \N__42553\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42548\,
            I => \N__42543\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42547\,
            I => \N__42540\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42537\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__42543\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42540\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__42537\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9350\ : CascadeMux
    port map (
            O => \N__42530\,
            I => \N__42527\
        );

    \I__9349\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42524\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__42524\,
            I => \N__42521\
        );

    \I__9347\ : Span4Mux_h
    port map (
            O => \N__42521\,
            I => \N__42518\
        );

    \I__9346\ : Odrv4
    port map (
            O => \N__42518\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__9345\ : CascadeMux
    port map (
            O => \N__42515\,
            I => \N__42511\
        );

    \I__9344\ : InMux
    port map (
            O => \N__42514\,
            I => \N__42507\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42511\,
            I => \N__42502\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42510\,
            I => \N__42502\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__42507\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__42502\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42497\,
            I => \N__42494\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__42494\,
            I => \N__42491\
        );

    \I__9337\ : Span4Mux_h
    port map (
            O => \N__42491\,
            I => \N__42488\
        );

    \I__9336\ : Odrv4
    port map (
            O => \N__42488\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42485\,
            I => \N__42482\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__42482\,
            I => \N__42479\
        );

    \I__9333\ : Odrv4
    port map (
            O => \N__42479\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__9332\ : CascadeMux
    port map (
            O => \N__42476\,
            I => \N__42462\
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__42475\,
            I => \N__42456\
        );

    \I__9330\ : CascadeMux
    port map (
            O => \N__42474\,
            I => \N__42453\
        );

    \I__9329\ : CascadeMux
    port map (
            O => \N__42473\,
            I => \N__42448\
        );

    \I__9328\ : CascadeMux
    port map (
            O => \N__42472\,
            I => \N__42434\
        );

    \I__9327\ : CascadeMux
    port map (
            O => \N__42471\,
            I => \N__42428\
        );

    \I__9326\ : CascadeMux
    port map (
            O => \N__42470\,
            I => \N__42425\
        );

    \I__9325\ : CascadeMux
    port map (
            O => \N__42469\,
            I => \N__42417\
        );

    \I__9324\ : CascadeMux
    port map (
            O => \N__42468\,
            I => \N__42413\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__42467\,
            I => \N__42408\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__42466\,
            I => \N__42404\
        );

    \I__9321\ : CascadeMux
    port map (
            O => \N__42465\,
            I => \N__42400\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42384\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42461\,
            I => \N__42373\
        );

    \I__9318\ : InMux
    port map (
            O => \N__42460\,
            I => \N__42373\
        );

    \I__9317\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42373\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42373\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42373\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42452\,
            I => \N__42370\
        );

    \I__9313\ : InMux
    port map (
            O => \N__42451\,
            I => \N__42359\
        );

    \I__9312\ : InMux
    port map (
            O => \N__42448\,
            I => \N__42359\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42447\,
            I => \N__42359\
        );

    \I__9310\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42359\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42359\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42342\
        );

    \I__9307\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42342\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42442\,
            I => \N__42342\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42342\
        );

    \I__9304\ : InMux
    port map (
            O => \N__42440\,
            I => \N__42342\
        );

    \I__9303\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42342\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42342\
        );

    \I__9301\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42342\
        );

    \I__9300\ : InMux
    port map (
            O => \N__42434\,
            I => \N__42339\
        );

    \I__9299\ : InMux
    port map (
            O => \N__42433\,
            I => \N__42328\
        );

    \I__9298\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42328\
        );

    \I__9297\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42328\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42328\
        );

    \I__9295\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42328\
        );

    \I__9294\ : CascadeMux
    port map (
            O => \N__42424\,
            I => \N__42315\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__42423\,
            I => \N__42311\
        );

    \I__9292\ : CascadeMux
    port map (
            O => \N__42422\,
            I => \N__42307\
        );

    \I__9291\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42291\
        );

    \I__9290\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42291\
        );

    \I__9289\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42274\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42274\
        );

    \I__9287\ : InMux
    port map (
            O => \N__42413\,
            I => \N__42274\
        );

    \I__9286\ : InMux
    port map (
            O => \N__42412\,
            I => \N__42274\
        );

    \I__9285\ : InMux
    port map (
            O => \N__42411\,
            I => \N__42274\
        );

    \I__9284\ : InMux
    port map (
            O => \N__42408\,
            I => \N__42274\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42407\,
            I => \N__42274\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42274\
        );

    \I__9281\ : InMux
    port map (
            O => \N__42403\,
            I => \N__42265\
        );

    \I__9280\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42265\
        );

    \I__9279\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42265\
        );

    \I__9278\ : InMux
    port map (
            O => \N__42398\,
            I => \N__42265\
        );

    \I__9277\ : CascadeMux
    port map (
            O => \N__42397\,
            I => \N__42262\
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__42396\,
            I => \N__42258\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__42395\,
            I => \N__42254\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__42394\,
            I => \N__42250\
        );

    \I__9273\ : CascadeMux
    port map (
            O => \N__42393\,
            I => \N__42238\
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__42392\,
            I => \N__42234\
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__42391\,
            I => \N__42230\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__42390\,
            I => \N__42226\
        );

    \I__9269\ : CascadeMux
    port map (
            O => \N__42389\,
            I => \N__42222\
        );

    \I__9268\ : CascadeMux
    port map (
            O => \N__42388\,
            I => \N__42218\
        );

    \I__9267\ : CascadeMux
    port map (
            O => \N__42387\,
            I => \N__42214\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__42384\,
            I => \N__42208\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__42373\,
            I => \N__42208\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__42370\,
            I => \N__42205\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__42359\,
            I => \N__42200\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__42342\,
            I => \N__42200\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__42339\,
            I => \N__42195\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42328\,
            I => \N__42195\
        );

    \I__9259\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42188\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42188\
        );

    \I__9257\ : InMux
    port map (
            O => \N__42325\,
            I => \N__42188\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__42324\,
            I => \N__42185\
        );

    \I__9255\ : CascadeMux
    port map (
            O => \N__42323\,
            I => \N__42179\
        );

    \I__9254\ : CascadeMux
    port map (
            O => \N__42322\,
            I => \N__42176\
        );

    \I__9253\ : CascadeMux
    port map (
            O => \N__42321\,
            I => \N__42173\
        );

    \I__9252\ : CascadeMux
    port map (
            O => \N__42320\,
            I => \N__42170\
        );

    \I__9251\ : CascadeMux
    port map (
            O => \N__42319\,
            I => \N__42167\
        );

    \I__9250\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42145\
        );

    \I__9249\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42145\
        );

    \I__9248\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42145\
        );

    \I__9247\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42145\
        );

    \I__9246\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42145\
        );

    \I__9245\ : InMux
    port map (
            O => \N__42307\,
            I => \N__42145\
        );

    \I__9244\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42145\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__42305\,
            I => \N__42140\
        );

    \I__9242\ : CascadeMux
    port map (
            O => \N__42304\,
            I => \N__42136\
        );

    \I__9241\ : CascadeMux
    port map (
            O => \N__42303\,
            I => \N__42132\
        );

    \I__9240\ : CascadeMux
    port map (
            O => \N__42302\,
            I => \N__42128\
        );

    \I__9239\ : CascadeMux
    port map (
            O => \N__42301\,
            I => \N__42124\
        );

    \I__9238\ : CascadeMux
    port map (
            O => \N__42300\,
            I => \N__42120\
        );

    \I__9237\ : CascadeMux
    port map (
            O => \N__42299\,
            I => \N__42116\
        );

    \I__9236\ : CascadeMux
    port map (
            O => \N__42298\,
            I => \N__42112\
        );

    \I__9235\ : CascadeMux
    port map (
            O => \N__42297\,
            I => \N__42108\
        );

    \I__9234\ : CascadeMux
    port map (
            O => \N__42296\,
            I => \N__42104\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__42291\,
            I => \N__42096\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__42274\,
            I => \N__42096\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__42265\,
            I => \N__42096\
        );

    \I__9230\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42079\
        );

    \I__9229\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42079\
        );

    \I__9228\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42079\
        );

    \I__9227\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42079\
        );

    \I__9226\ : InMux
    port map (
            O => \N__42254\,
            I => \N__42079\
        );

    \I__9225\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42079\
        );

    \I__9224\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42079\
        );

    \I__9223\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42079\
        );

    \I__9222\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42070\
        );

    \I__9221\ : InMux
    port map (
            O => \N__42247\,
            I => \N__42070\
        );

    \I__9220\ : InMux
    port map (
            O => \N__42246\,
            I => \N__42070\
        );

    \I__9219\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42070\
        );

    \I__9218\ : InMux
    port map (
            O => \N__42244\,
            I => \N__42061\
        );

    \I__9217\ : InMux
    port map (
            O => \N__42243\,
            I => \N__42061\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42061\
        );

    \I__9215\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42061\
        );

    \I__9214\ : InMux
    port map (
            O => \N__42238\,
            I => \N__42044\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42237\,
            I => \N__42044\
        );

    \I__9212\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42044\
        );

    \I__9211\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42044\
        );

    \I__9210\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42044\
        );

    \I__9209\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42044\
        );

    \I__9208\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42044\
        );

    \I__9207\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42044\
        );

    \I__9206\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42031\
        );

    \I__9205\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42031\
        );

    \I__9204\ : InMux
    port map (
            O => \N__42218\,
            I => \N__42031\
        );

    \I__9203\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42031\
        );

    \I__9202\ : InMux
    port map (
            O => \N__42214\,
            I => \N__42031\
        );

    \I__9201\ : InMux
    port map (
            O => \N__42213\,
            I => \N__42031\
        );

    \I__9200\ : Span12Mux_s11_h
    port map (
            O => \N__42208\,
            I => \N__42028\
        );

    \I__9199\ : Span4Mux_v
    port map (
            O => \N__42205\,
            I => \N__42019\
        );

    \I__9198\ : Span4Mux_h
    port map (
            O => \N__42200\,
            I => \N__42019\
        );

    \I__9197\ : Span4Mux_v
    port map (
            O => \N__42195\,
            I => \N__42019\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__42188\,
            I => \N__42019\
        );

    \I__9195\ : InMux
    port map (
            O => \N__42185\,
            I => \N__42010\
        );

    \I__9194\ : InMux
    port map (
            O => \N__42184\,
            I => \N__42010\
        );

    \I__9193\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42010\
        );

    \I__9192\ : InMux
    port map (
            O => \N__42182\,
            I => \N__42010\
        );

    \I__9191\ : InMux
    port map (
            O => \N__42179\,
            I => \N__42003\
        );

    \I__9190\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42003\
        );

    \I__9189\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42003\
        );

    \I__9188\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42000\
        );

    \I__9187\ : InMux
    port map (
            O => \N__42167\,
            I => \N__41985\
        );

    \I__9186\ : InMux
    port map (
            O => \N__42166\,
            I => \N__41985\
        );

    \I__9185\ : InMux
    port map (
            O => \N__42165\,
            I => \N__41985\
        );

    \I__9184\ : InMux
    port map (
            O => \N__42164\,
            I => \N__41985\
        );

    \I__9183\ : InMux
    port map (
            O => \N__42163\,
            I => \N__41985\
        );

    \I__9182\ : InMux
    port map (
            O => \N__42162\,
            I => \N__41985\
        );

    \I__9181\ : InMux
    port map (
            O => \N__42161\,
            I => \N__41985\
        );

    \I__9180\ : InMux
    port map (
            O => \N__42160\,
            I => \N__41982\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__42145\,
            I => \N__41979\
        );

    \I__9178\ : InMux
    port map (
            O => \N__42144\,
            I => \N__41962\
        );

    \I__9177\ : InMux
    port map (
            O => \N__42143\,
            I => \N__41962\
        );

    \I__9176\ : InMux
    port map (
            O => \N__42140\,
            I => \N__41962\
        );

    \I__9175\ : InMux
    port map (
            O => \N__42139\,
            I => \N__41962\
        );

    \I__9174\ : InMux
    port map (
            O => \N__42136\,
            I => \N__41962\
        );

    \I__9173\ : InMux
    port map (
            O => \N__42135\,
            I => \N__41962\
        );

    \I__9172\ : InMux
    port map (
            O => \N__42132\,
            I => \N__41962\
        );

    \I__9171\ : InMux
    port map (
            O => \N__42131\,
            I => \N__41962\
        );

    \I__9170\ : InMux
    port map (
            O => \N__42128\,
            I => \N__41945\
        );

    \I__9169\ : InMux
    port map (
            O => \N__42127\,
            I => \N__41945\
        );

    \I__9168\ : InMux
    port map (
            O => \N__42124\,
            I => \N__41945\
        );

    \I__9167\ : InMux
    port map (
            O => \N__42123\,
            I => \N__41945\
        );

    \I__9166\ : InMux
    port map (
            O => \N__42120\,
            I => \N__41945\
        );

    \I__9165\ : InMux
    port map (
            O => \N__42119\,
            I => \N__41945\
        );

    \I__9164\ : InMux
    port map (
            O => \N__42116\,
            I => \N__41945\
        );

    \I__9163\ : InMux
    port map (
            O => \N__42115\,
            I => \N__41945\
        );

    \I__9162\ : InMux
    port map (
            O => \N__42112\,
            I => \N__41932\
        );

    \I__9161\ : InMux
    port map (
            O => \N__42111\,
            I => \N__41932\
        );

    \I__9160\ : InMux
    port map (
            O => \N__42108\,
            I => \N__41932\
        );

    \I__9159\ : InMux
    port map (
            O => \N__42107\,
            I => \N__41932\
        );

    \I__9158\ : InMux
    port map (
            O => \N__42104\,
            I => \N__41932\
        );

    \I__9157\ : InMux
    port map (
            O => \N__42103\,
            I => \N__41932\
        );

    \I__9156\ : Span12Mux_s11_h
    port map (
            O => \N__42096\,
            I => \N__41919\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__42079\,
            I => \N__41919\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__42070\,
            I => \N__41919\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__42061\,
            I => \N__41919\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__42044\,
            I => \N__41919\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__42031\,
            I => \N__41919\
        );

    \I__9150\ : Odrv12
    port map (
            O => \N__42028\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__42019\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__42010\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__42003\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__42000\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41985\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__41982\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__41979\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__41962\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__41945\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__41932\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9139\ : Odrv12
    port map (
            O => \N__41919\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__9138\ : CascadeMux
    port map (
            O => \N__41894\,
            I => \N__41891\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41888\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41888\,
            I => \N__41885\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__41885\,
            I => \N__41882\
        );

    \I__9134\ : Odrv4
    port map (
            O => \N__41882\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__41879\,
            I => \N__41875\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41878\,
            I => \N__41867\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41867\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41867\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__41867\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41849\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41840\
        );

    \I__9126\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41827\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41827\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41827\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41827\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41827\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41857\,
            I => \N__41827\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41856\,
            I => \N__41816\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41855\,
            I => \N__41816\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41816\
        );

    \I__9117\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41816\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41816\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41849\,
            I => \N__41813\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41848\,
            I => \N__41808\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41847\,
            I => \N__41808\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41793\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41845\,
            I => \N__41793\
        );

    \I__9110\ : InMux
    port map (
            O => \N__41844\,
            I => \N__41793\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41793\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__41840\,
            I => \N__41786\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__41827\,
            I => \N__41786\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__41816\,
            I => \N__41786\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__41813\,
            I => \N__41781\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__41808\,
            I => \N__41781\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41778\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41767\
        );

    \I__9101\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41767\
        );

    \I__9100\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41767\
        );

    \I__9099\ : InMux
    port map (
            O => \N__41803\,
            I => \N__41767\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41802\,
            I => \N__41767\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41760\
        );

    \I__9096\ : Span4Mux_v
    port map (
            O => \N__41786\,
            I => \N__41760\
        );

    \I__9095\ : Span4Mux_h
    port map (
            O => \N__41781\,
            I => \N__41760\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41778\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__41767\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__41760\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41750\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__41750\,
            I => \N__41745\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41742\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41748\,
            I => \N__41739\
        );

    \I__9087\ : Odrv4
    port map (
            O => \N__41745\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41742\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__41739\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41732\,
            I => \N__41729\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__41729\,
            I => \N__41724\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41728\,
            I => \N__41721\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41727\,
            I => \N__41718\
        );

    \I__9080\ : Odrv4
    port map (
            O => \N__41724\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__41721\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41718\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41711\,
            I => \N__41708\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__41708\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__9075\ : CascadeMux
    port map (
            O => \N__41705\,
            I => \N__41702\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41702\,
            I => \N__41699\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__41699\,
            I => \N__41695\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41691\
        );

    \I__9071\ : Span4Mux_h
    port map (
            O => \N__41695\,
            I => \N__41688\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41694\,
            I => \N__41685\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__41691\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9068\ : Odrv4
    port map (
            O => \N__41688\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__41685\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41678\,
            I => \N__41673\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41677\,
            I => \N__41670\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41676\,
            I => \N__41667\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__41673\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__41670\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41667\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__41660\,
            I => \N__41657\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41654\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41654\,
            I => \N__41650\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41647\
        );

    \I__9056\ : Span4Mux_v
    port map (
            O => \N__41650\,
            I => \N__41641\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41647\,
            I => \N__41641\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41638\
        );

    \I__9053\ : Odrv4
    port map (
            O => \N__41641\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41638\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9051\ : InMux
    port map (
            O => \N__41633\,
            I => \N__41630\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__41630\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41627\,
            I => \N__41624\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__41624\,
            I => \N__41619\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41623\,
            I => \N__41616\
        );

    \I__9046\ : InMux
    port map (
            O => \N__41622\,
            I => \N__41613\
        );

    \I__9045\ : Odrv12
    port map (
            O => \N__41619\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__41616\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__41613\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41603\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__41603\,
            I => \N__41599\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41595\
        );

    \I__9039\ : Span4Mux_h
    port map (
            O => \N__41599\,
            I => \N__41592\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41589\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41595\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__41592\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__41589\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__41582\,
            I => \N__41579\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41576\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__41576\,
            I => \N__41573\
        );

    \I__9031\ : Span4Mux_v
    port map (
            O => \N__41573\,
            I => \N__41569\
        );

    \I__9030\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41566\
        );

    \I__9029\ : Span4Mux_h
    port map (
            O => \N__41569\,
            I => \N__41562\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__41566\,
            I => \N__41559\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41556\
        );

    \I__9026\ : Odrv4
    port map (
            O => \N__41562\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9025\ : Odrv4
    port map (
            O => \N__41559\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__41556\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9023\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41546\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__41546\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__9021\ : CascadeMux
    port map (
            O => \N__41543\,
            I => \N__41539\
        );

    \I__9020\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41536\
        );

    \I__9019\ : InMux
    port map (
            O => \N__41539\,
            I => \N__41533\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__41536\,
            I => \N__41529\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__41533\,
            I => \N__41526\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41532\,
            I => \N__41523\
        );

    \I__9015\ : Odrv4
    port map (
            O => \N__41529\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__41526\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41523\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9012\ : InMux
    port map (
            O => \N__41516\,
            I => \N__41512\
        );

    \I__9011\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41509\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__41512\,
            I => \N__41503\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__41509\,
            I => \N__41503\
        );

    \I__9008\ : InMux
    port map (
            O => \N__41508\,
            I => \N__41500\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__41503\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__41500\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9005\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41492\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__41492\,
            I => \N__41487\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41484\
        );

    \I__9002\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41481\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__41487\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41484\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41481\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41471\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__41471\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__8996\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41464\
        );

    \I__8995\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41461\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__41464\,
            I => \N__41457\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__41461\,
            I => \N__41454\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41460\,
            I => \N__41451\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__41457\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__41454\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__41451\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8988\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41441\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__41441\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41438\,
            I => \N__41435\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__41435\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__41432\,
            I => \N__41429\
        );

    \I__8983\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41426\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__41426\,
            I => \N__41421\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41425\,
            I => \N__41416\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41416\
        );

    \I__8979\ : Odrv4
    port map (
            O => \N__41421\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__41416\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8977\ : CascadeMux
    port map (
            O => \N__41411\,
            I => \N__41408\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41408\,
            I => \N__41404\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41407\,
            I => \N__41401\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41404\,
            I => \N__41397\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__41401\,
            I => \N__41394\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41400\,
            I => \N__41391\
        );

    \I__8971\ : Odrv12
    port map (
            O => \N__41397\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8970\ : Odrv4
    port map (
            O => \N__41394\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41391\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41381\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__41381\,
            I => \N__41376\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41373\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41370\
        );

    \I__8964\ : Odrv4
    port map (
            O => \N__41376\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__41373\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__41370\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__8961\ : InMux
    port map (
            O => \N__41363\,
            I => \N__41359\
        );

    \I__8960\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41356\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__41359\,
            I => \N__41353\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__41356\,
            I => \N__41348\
        );

    \I__8957\ : Span4Mux_h
    port map (
            O => \N__41353\,
            I => \N__41345\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41352\,
            I => \N__41340\
        );

    \I__8955\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41340\
        );

    \I__8954\ : Odrv12
    port map (
            O => \N__41348\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__41345\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41340\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41329\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41326\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__41329\,
            I => \N__41322\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__41326\,
            I => \N__41319\
        );

    \I__8947\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41316\
        );

    \I__8946\ : Odrv4
    port map (
            O => \N__41322\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8945\ : Odrv4
    port map (
            O => \N__41319\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__41316\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41309\,
            I => \N__41305\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41308\,
            I => \N__41302\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__41305\,
            I => \N__41298\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__41302\,
            I => \N__41295\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41292\
        );

    \I__8938\ : Odrv4
    port map (
            O => \N__41298\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__41295\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__41292\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__8935\ : InMux
    port map (
            O => \N__41285\,
            I => \N__41280\
        );

    \I__8934\ : CascadeMux
    port map (
            O => \N__41284\,
            I => \N__41277\
        );

    \I__8933\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41273\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__41280\,
            I => \N__41270\
        );

    \I__8931\ : InMux
    port map (
            O => \N__41277\,
            I => \N__41267\
        );

    \I__8930\ : InMux
    port map (
            O => \N__41276\,
            I => \N__41263\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__41273\,
            I => \N__41260\
        );

    \I__8928\ : Span4Mux_v
    port map (
            O => \N__41270\,
            I => \N__41257\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__41267\,
            I => \N__41254\
        );

    \I__8926\ : InMux
    port map (
            O => \N__41266\,
            I => \N__41251\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__41263\,
            I => \N__41248\
        );

    \I__8924\ : Span4Mux_v
    port map (
            O => \N__41260\,
            I => \N__41245\
        );

    \I__8923\ : Span4Mux_h
    port map (
            O => \N__41257\,
            I => \N__41242\
        );

    \I__8922\ : Span4Mux_h
    port map (
            O => \N__41254\,
            I => \N__41237\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__41251\,
            I => \N__41237\
        );

    \I__8920\ : Span4Mux_v
    port map (
            O => \N__41248\,
            I => \N__41230\
        );

    \I__8919\ : Span4Mux_h
    port map (
            O => \N__41245\,
            I => \N__41230\
        );

    \I__8918\ : Span4Mux_h
    port map (
            O => \N__41242\,
            I => \N__41230\
        );

    \I__8917\ : Odrv4
    port map (
            O => \N__41237\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8916\ : Odrv4
    port map (
            O => \N__41230\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41225\,
            I => \N__41222\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__41222\,
            I => \N__41219\
        );

    \I__8913\ : Span4Mux_v
    port map (
            O => \N__41219\,
            I => \N__41216\
        );

    \I__8912\ : Sp12to4
    port map (
            O => \N__41216\,
            I => \N__41213\
        );

    \I__8911\ : Span12Mux_h
    port map (
            O => \N__41213\,
            I => \N__41210\
        );

    \I__8910\ : Odrv12
    port map (
            O => \N__41210\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__8909\ : CascadeMux
    port map (
            O => \N__41207\,
            I => \N__41204\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41200\
        );

    \I__8907\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41196\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__41200\,
            I => \N__41193\
        );

    \I__8905\ : InMux
    port map (
            O => \N__41199\,
            I => \N__41190\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__41196\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8903\ : Odrv4
    port map (
            O => \N__41193\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__41190\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8901\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41176\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41176\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41173\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__41176\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__41173\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8896\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41164\
        );

    \I__8895\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41161\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41164\,
            I => \N__41157\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41161\,
            I => \N__41154\
        );

    \I__8892\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41151\
        );

    \I__8891\ : Odrv4
    port map (
            O => \N__41157\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8890\ : Odrv12
    port map (
            O => \N__41154\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__41151\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8888\ : InMux
    port map (
            O => \N__41144\,
            I => \N__41141\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__41141\,
            I => \N__41137\
        );

    \I__8886\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41134\
        );

    \I__8885\ : Span4Mux_h
    port map (
            O => \N__41137\,
            I => \N__41131\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__41134\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__41131\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8882\ : CascadeMux
    port map (
            O => \N__41126\,
            I => \N__41123\
        );

    \I__8881\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41118\
        );

    \I__8880\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41115\
        );

    \I__8879\ : InMux
    port map (
            O => \N__41121\,
            I => \N__41112\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__41118\,
            I => \N__41107\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__41115\,
            I => \N__41107\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__41112\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__41107\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8874\ : InMux
    port map (
            O => \N__41102\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8873\ : InMux
    port map (
            O => \N__41099\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8872\ : CEMux
    port map (
            O => \N__41096\,
            I => \N__41091\
        );

    \I__8871\ : CEMux
    port map (
            O => \N__41095\,
            I => \N__41088\
        );

    \I__8870\ : CEMux
    port map (
            O => \N__41094\,
            I => \N__41084\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__41091\,
            I => \N__41080\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__41088\,
            I => \N__41077\
        );

    \I__8867\ : CEMux
    port map (
            O => \N__41087\,
            I => \N__41074\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__41084\,
            I => \N__41071\
        );

    \I__8865\ : CEMux
    port map (
            O => \N__41083\,
            I => \N__41068\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__41080\,
            I => \N__41061\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__41077\,
            I => \N__41061\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__41074\,
            I => \N__41061\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__41071\,
            I => \N__41058\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__41068\,
            I => \N__41055\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__41061\,
            I => \N__41052\
        );

    \I__8858\ : Span4Mux_v
    port map (
            O => \N__41058\,
            I => \N__41049\
        );

    \I__8857\ : Span4Mux_v
    port map (
            O => \N__41055\,
            I => \N__41046\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__41052\,
            I => \N__41043\
        );

    \I__8855\ : Odrv4
    port map (
            O => \N__41049\,
            I => \delay_measurement_inst.delay_hc_timer.N_201_i\
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__41046\,
            I => \delay_measurement_inst.delay_hc_timer.N_201_i\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__41043\,
            I => \delay_measurement_inst.delay_hc_timer.N_201_i\
        );

    \I__8852\ : InMux
    port map (
            O => \N__41036\,
            I => \N__41030\
        );

    \I__8851\ : InMux
    port map (
            O => \N__41035\,
            I => \N__41030\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__41030\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__8849\ : InMux
    port map (
            O => \N__41027\,
            I => \N__41024\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__41024\,
            I => \N__41020\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41023\,
            I => \N__41017\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__41020\,
            I => \N__41011\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__41017\,
            I => \N__41011\
        );

    \I__8844\ : InMux
    port map (
            O => \N__41016\,
            I => \N__41008\
        );

    \I__8843\ : Span4Mux_v
    port map (
            O => \N__41011\,
            I => \N__41002\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__41008\,
            I => \N__41002\
        );

    \I__8841\ : InMux
    port map (
            O => \N__41007\,
            I => \N__40999\
        );

    \I__8840\ : Span4Mux_h
    port map (
            O => \N__41002\,
            I => \N__40996\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__40999\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__40996\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8837\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40987\
        );

    \I__8836\ : InMux
    port map (
            O => \N__40990\,
            I => \N__40983\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40987\,
            I => \N__40980\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40986\,
            I => \N__40977\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40983\,
            I => \N__40974\
        );

    \I__8832\ : Span4Mux_v
    port map (
            O => \N__40980\,
            I => \N__40971\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40977\,
            I => \N__40966\
        );

    \I__8830\ : Span4Mux_v
    port map (
            O => \N__40974\,
            I => \N__40966\
        );

    \I__8829\ : Odrv4
    port map (
            O => \N__40971\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8828\ : Odrv4
    port map (
            O => \N__40966\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40956\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40960\,
            I => \N__40953\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40950\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40956\,
            I => \N__40945\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40953\,
            I => \N__40945\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__40950\,
            I => \N__40942\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__40945\,
            I => \N__40939\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__40942\,
            I => \N__40936\
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__40939\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__8818\ : Odrv4
    port map (
            O => \N__40936\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__8817\ : CascadeMux
    port map (
            O => \N__40931\,
            I => \N__40927\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40930\,
            I => \N__40922\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40927\,
            I => \N__40922\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40922\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40919\,
            I => \N__40916\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__40916\,
            I => \N__40912\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40915\,
            I => \N__40909\
        );

    \I__8810\ : Span4Mux_v
    port map (
            O => \N__40912\,
            I => \N__40905\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__40909\,
            I => \N__40902\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40908\,
            I => \N__40899\
        );

    \I__8807\ : Span4Mux_h
    port map (
            O => \N__40905\,
            I => \N__40894\
        );

    \I__8806\ : Span4Mux_h
    port map (
            O => \N__40902\,
            I => \N__40894\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__40899\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__8804\ : Odrv4
    port map (
            O => \N__40894\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40889\,
            I => \N__40884\
        );

    \I__8802\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40881\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40878\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__40884\,
            I => \N__40875\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__40881\,
            I => \N__40868\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__40878\,
            I => \N__40868\
        );

    \I__8797\ : Span4Mux_h
    port map (
            O => \N__40875\,
            I => \N__40868\
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__40868\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40859\
        );

    \I__8794\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40859\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40859\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__8792\ : CascadeMux
    port map (
            O => \N__40856\,
            I => \N__40853\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40853\,
            I => \N__40850\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__40850\,
            I => \N__40847\
        );

    \I__8789\ : Odrv4
    port map (
            O => \N__40847\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40841\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__40841\,
            I => \N__40838\
        );

    \I__8786\ : Span4Mux_h
    port map (
            O => \N__40838\,
            I => \N__40835\
        );

    \I__8785\ : Odrv4
    port map (
            O => \N__40835\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__8784\ : CascadeMux
    port map (
            O => \N__40832\,
            I => \N__40829\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40829\,
            I => \N__40824\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40828\,
            I => \N__40821\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40827\,
            I => \N__40818\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40824\,
            I => \N__40813\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40821\,
            I => \N__40813\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40818\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8777\ : Odrv4
    port map (
            O => \N__40813\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40808\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40805\,
            I => \N__40798\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40798\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40795\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__40798\,
            I => \N__40792\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40795\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8770\ : Odrv4
    port map (
            O => \N__40792\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40787\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40778\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40778\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__40778\,
            I => \N__40774\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40771\
        );

    \I__8764\ : Span4Mux_h
    port map (
            O => \N__40774\,
            I => \N__40768\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40771\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8762\ : Odrv4
    port map (
            O => \N__40768\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40763\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__40760\,
            I => \N__40756\
        );

    \I__8759\ : CascadeMux
    port map (
            O => \N__40759\,
            I => \N__40753\
        );

    \I__8758\ : InMux
    port map (
            O => \N__40756\,
            I => \N__40748\
        );

    \I__8757\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40748\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40748\,
            I => \N__40744\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40741\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__40744\,
            I => \N__40738\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40741\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8752\ : Odrv4
    port map (
            O => \N__40738\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40733\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8750\ : CascadeMux
    port map (
            O => \N__40730\,
            I => \N__40726\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__40729\,
            I => \N__40723\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40726\,
            I => \N__40718\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40723\,
            I => \N__40718\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__40718\,
            I => \N__40714\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40711\
        );

    \I__8744\ : Span4Mux_v
    port map (
            O => \N__40714\,
            I => \N__40708\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40711\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__40708\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40703\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8740\ : CascadeMux
    port map (
            O => \N__40700\,
            I => \N__40697\
        );

    \I__8739\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40694\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__40694\,
            I => \N__40689\
        );

    \I__8737\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40686\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40683\
        );

    \I__8735\ : Span4Mux_v
    port map (
            O => \N__40689\,
            I => \N__40678\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40686\,
            I => \N__40678\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40683\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__40678\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8731\ : InMux
    port map (
            O => \N__40673\,
            I => \bfn_16_23_0_\
        );

    \I__8730\ : CascadeMux
    port map (
            O => \N__40670\,
            I => \N__40667\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40664\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40664\,
            I => \N__40659\
        );

    \I__8727\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40656\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40662\,
            I => \N__40653\
        );

    \I__8725\ : Span4Mux_v
    port map (
            O => \N__40659\,
            I => \N__40648\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__40656\,
            I => \N__40648\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40653\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8722\ : Odrv4
    port map (
            O => \N__40648\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40643\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40640\,
            I => \N__40636\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40633\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__40636\,
            I => \N__40630\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__40633\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8716\ : Odrv4
    port map (
            O => \N__40630\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8715\ : CascadeMux
    port map (
            O => \N__40625\,
            I => \N__40622\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40617\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40614\
        );

    \I__8712\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40611\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40617\,
            I => \N__40606\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__40614\,
            I => \N__40606\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__40611\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__40606\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40601\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8706\ : InMux
    port map (
            O => \N__40598\,
            I => \N__40591\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40591\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40596\,
            I => \N__40588\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40591\,
            I => \N__40585\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40588\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__40585\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8700\ : InMux
    port map (
            O => \N__40580\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8699\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40570\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40570\
        );

    \I__8697\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40567\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__40570\,
            I => \N__40564\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__40567\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8694\ : Odrv4
    port map (
            O => \N__40564\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40559\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8692\ : CascadeMux
    port map (
            O => \N__40556\,
            I => \N__40552\
        );

    \I__8691\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40548\
        );

    \I__8690\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40545\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40542\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__40548\,
            I => \N__40537\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__40545\,
            I => \N__40537\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40542\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__40537\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8684\ : InMux
    port map (
            O => \N__40532\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__40529\,
            I => \N__40525\
        );

    \I__8682\ : InMux
    port map (
            O => \N__40528\,
            I => \N__40521\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40518\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40515\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__40521\,
            I => \N__40510\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40518\,
            I => \N__40510\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__40515\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8676\ : Odrv4
    port map (
            O => \N__40510\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8675\ : InMux
    port map (
            O => \N__40505\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__40502\,
            I => \N__40498\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__40501\,
            I => \N__40495\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40498\,
            I => \N__40489\
        );

    \I__8671\ : InMux
    port map (
            O => \N__40495\,
            I => \N__40489\
        );

    \I__8670\ : InMux
    port map (
            O => \N__40494\,
            I => \N__40486\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__40489\,
            I => \N__40483\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__40486\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__40483\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8666\ : InMux
    port map (
            O => \N__40478\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8665\ : CascadeMux
    port map (
            O => \N__40475\,
            I => \N__40471\
        );

    \I__8664\ : CascadeMux
    port map (
            O => \N__40474\,
            I => \N__40468\
        );

    \I__8663\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40462\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40468\,
            I => \N__40462\
        );

    \I__8661\ : InMux
    port map (
            O => \N__40467\,
            I => \N__40459\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__40462\,
            I => \N__40456\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__40459\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8658\ : Odrv4
    port map (
            O => \N__40456\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8657\ : InMux
    port map (
            O => \N__40451\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__40448\,
            I => \N__40445\
        );

    \I__8655\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40442\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40442\,
            I => \N__40437\
        );

    \I__8653\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40434\
        );

    \I__8652\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40431\
        );

    \I__8651\ : Span4Mux_v
    port map (
            O => \N__40437\,
            I => \N__40426\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__40434\,
            I => \N__40426\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__40431\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8648\ : Odrv4
    port map (
            O => \N__40426\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8647\ : InMux
    port map (
            O => \N__40421\,
            I => \bfn_16_22_0_\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__40418\,
            I => \N__40415\
        );

    \I__8645\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40411\
        );

    \I__8644\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40408\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__40411\,
            I => \N__40404\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__40408\,
            I => \N__40401\
        );

    \I__8641\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40398\
        );

    \I__8640\ : Span4Mux_v
    port map (
            O => \N__40404\,
            I => \N__40395\
        );

    \I__8639\ : Span4Mux_h
    port map (
            O => \N__40401\,
            I => \N__40392\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__40398\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8637\ : Odrv4
    port map (
            O => \N__40395\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__40392\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8635\ : InMux
    port map (
            O => \N__40385\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8634\ : CascadeMux
    port map (
            O => \N__40382\,
            I => \N__40379\
        );

    \I__8633\ : InMux
    port map (
            O => \N__40379\,
            I => \N__40374\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40371\
        );

    \I__8631\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40368\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__40374\,
            I => \N__40363\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__40371\,
            I => \N__40363\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__40368\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8627\ : Odrv4
    port map (
            O => \N__40363\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40358\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40355\,
            I => \N__40348\
        );

    \I__8624\ : InMux
    port map (
            O => \N__40354\,
            I => \N__40348\
        );

    \I__8623\ : InMux
    port map (
            O => \N__40353\,
            I => \N__40345\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__40348\,
            I => \N__40342\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__40345\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__40342\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8619\ : InMux
    port map (
            O => \N__40337\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__40334\,
            I => \N__40330\
        );

    \I__8617\ : CascadeMux
    port map (
            O => \N__40333\,
            I => \N__40327\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40330\,
            I => \N__40322\
        );

    \I__8615\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40322\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__40322\,
            I => \N__40318\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40321\,
            I => \N__40315\
        );

    \I__8612\ : Span4Mux_v
    port map (
            O => \N__40318\,
            I => \N__40312\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__40315\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8610\ : Odrv4
    port map (
            O => \N__40312\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40307\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8608\ : CascadeMux
    port map (
            O => \N__40304\,
            I => \N__40300\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40303\,
            I => \N__40296\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40293\
        );

    \I__8605\ : InMux
    port map (
            O => \N__40299\,
            I => \N__40290\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__40296\,
            I => \N__40285\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40293\,
            I => \N__40285\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__40290\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__40285\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8600\ : InMux
    port map (
            O => \N__40280\,
            I => \N__40274\
        );

    \I__8599\ : InMux
    port map (
            O => \N__40279\,
            I => \N__40271\
        );

    \I__8598\ : InMux
    port map (
            O => \N__40278\,
            I => \N__40268\
        );

    \I__8597\ : InMux
    port map (
            O => \N__40277\,
            I => \N__40265\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__40274\,
            I => \N__40262\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40271\,
            I => \N__40259\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__40268\,
            I => \N__40256\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__40265\,
            I => \N__40253\
        );

    \I__8592\ : Span4Mux_v
    port map (
            O => \N__40262\,
            I => \N__40250\
        );

    \I__8591\ : Span4Mux_h
    port map (
            O => \N__40259\,
            I => \N__40247\
        );

    \I__8590\ : Span4Mux_h
    port map (
            O => \N__40256\,
            I => \N__40244\
        );

    \I__8589\ : Odrv12
    port map (
            O => \N__40253\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__8588\ : Odrv4
    port map (
            O => \N__40250\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__40247\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__8586\ : Odrv4
    port map (
            O => \N__40244\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__8585\ : InMux
    port map (
            O => \N__40235\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40225\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40231\,
            I => \N__40225\
        );

    \I__8582\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40222\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40225\,
            I => \N__40219\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__40222\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__40219\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8578\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40208\
        );

    \I__8577\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40205\
        );

    \I__8576\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40202\
        );

    \I__8575\ : InMux
    port map (
            O => \N__40211\,
            I => \N__40199\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__40208\,
            I => \N__40196\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__40205\,
            I => \N__40191\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__40202\,
            I => \N__40191\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40188\
        );

    \I__8570\ : Span12Mux_h
    port map (
            O => \N__40196\,
            I => \N__40185\
        );

    \I__8569\ : Span4Mux_v
    port map (
            O => \N__40191\,
            I => \N__40182\
        );

    \I__8568\ : Span4Mux_h
    port map (
            O => \N__40188\,
            I => \N__40179\
        );

    \I__8567\ : Odrv12
    port map (
            O => \N__40185\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__40182\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__40179\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8564\ : InMux
    port map (
            O => \N__40172\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__40169\,
            I => \N__40165\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__40168\,
            I => \N__40162\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40165\,
            I => \N__40156\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40162\,
            I => \N__40156\
        );

    \I__8559\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40153\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__40156\,
            I => \N__40150\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__40153\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__8556\ : Odrv4
    port map (
            O => \N__40150\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__8555\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40141\
        );

    \I__8554\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40136\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__40141\,
            I => \N__40133\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40130\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40127\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40136\,
            I => \N__40124\
        );

    \I__8549\ : Span4Mux_v
    port map (
            O => \N__40133\,
            I => \N__40119\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__40130\,
            I => \N__40119\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__40127\,
            I => \N__40116\
        );

    \I__8546\ : Span4Mux_h
    port map (
            O => \N__40124\,
            I => \N__40111\
        );

    \I__8545\ : Span4Mux_h
    port map (
            O => \N__40119\,
            I => \N__40111\
        );

    \I__8544\ : Span4Mux_h
    port map (
            O => \N__40116\,
            I => \N__40108\
        );

    \I__8543\ : Odrv4
    port map (
            O => \N__40111\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__8542\ : Odrv4
    port map (
            O => \N__40108\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__8541\ : InMux
    port map (
            O => \N__40103\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__40100\,
            I => \N__40096\
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__40099\,
            I => \N__40093\
        );

    \I__8538\ : InMux
    port map (
            O => \N__40096\,
            I => \N__40087\
        );

    \I__8537\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40087\
        );

    \I__8536\ : InMux
    port map (
            O => \N__40092\,
            I => \N__40084\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__40087\,
            I => \N__40081\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40084\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__8533\ : Odrv4
    port map (
            O => \N__40081\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__8532\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40071\
        );

    \I__8531\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40067\
        );

    \I__8530\ : InMux
    port map (
            O => \N__40074\,
            I => \N__40064\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__40071\,
            I => \N__40061\
        );

    \I__8528\ : InMux
    port map (
            O => \N__40070\,
            I => \N__40058\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__40067\,
            I => \N__40055\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__40064\,
            I => \N__40052\
        );

    \I__8525\ : Span4Mux_v
    port map (
            O => \N__40061\,
            I => \N__40049\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__40058\,
            I => \N__40044\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__40055\,
            I => \N__40044\
        );

    \I__8522\ : Span4Mux_h
    port map (
            O => \N__40052\,
            I => \N__40041\
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__40049\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__40044\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__40041\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8518\ : InMux
    port map (
            O => \N__40034\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8517\ : CascadeMux
    port map (
            O => \N__40031\,
            I => \N__40028\
        );

    \I__8516\ : InMux
    port map (
            O => \N__40028\,
            I => \N__40025\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__40025\,
            I => \N__40020\
        );

    \I__8514\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40017\
        );

    \I__8513\ : InMux
    port map (
            O => \N__40023\,
            I => \N__40014\
        );

    \I__8512\ : Span4Mux_v
    port map (
            O => \N__40020\,
            I => \N__40009\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__40017\,
            I => \N__40009\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__40014\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__40009\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8508\ : InMux
    port map (
            O => \N__40004\,
            I => \N__39998\
        );

    \I__8507\ : InMux
    port map (
            O => \N__40003\,
            I => \N__39995\
        );

    \I__8506\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39992\
        );

    \I__8505\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39989\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39998\,
            I => \N__39986\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__39995\,
            I => \N__39983\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__39992\,
            I => \N__39980\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39989\,
            I => \N__39977\
        );

    \I__8500\ : Span4Mux_v
    port map (
            O => \N__39986\,
            I => \N__39972\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__39983\,
            I => \N__39972\
        );

    \I__8498\ : Span4Mux_h
    port map (
            O => \N__39980\,
            I => \N__39967\
        );

    \I__8497\ : Span4Mux_h
    port map (
            O => \N__39977\,
            I => \N__39967\
        );

    \I__8496\ : Odrv4
    port map (
            O => \N__39972\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__39967\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__8494\ : InMux
    port map (
            O => \N__39962\,
            I => \bfn_16_21_0_\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__39959\,
            I => \N__39956\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39956\,
            I => \N__39953\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39953\,
            I => \N__39948\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39952\,
            I => \N__39945\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39942\
        );

    \I__8488\ : Span4Mux_v
    port map (
            O => \N__39948\,
            I => \N__39937\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39945\,
            I => \N__39937\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__39942\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__39937\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39924\
        );

    \I__8482\ : InMux
    port map (
            O => \N__39928\,
            I => \N__39921\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39917\
        );

    \I__8480\ : Span4Mux_h
    port map (
            O => \N__39924\,
            I => \N__39912\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__39921\,
            I => \N__39912\
        );

    \I__8478\ : CascadeMux
    port map (
            O => \N__39920\,
            I => \N__39909\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39917\,
            I => \N__39906\
        );

    \I__8476\ : Span4Mux_h
    port map (
            O => \N__39912\,
            I => \N__39903\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39900\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__39906\,
            I => \N__39895\
        );

    \I__8473\ : Span4Mux_v
    port map (
            O => \N__39903\,
            I => \N__39895\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__39900\,
            I => \N__39892\
        );

    \I__8471\ : Span4Mux_v
    port map (
            O => \N__39895\,
            I => \N__39889\
        );

    \I__8470\ : Span4Mux_h
    port map (
            O => \N__39892\,
            I => \N__39886\
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__39889\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__39886\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39881\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8466\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39875\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39870\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39865\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39865\
        );

    \I__8462\ : Odrv4
    port map (
            O => \N__39870\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39865\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39857\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__39857\,
            I => \N__39853\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39856\,
            I => \N__39850\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__39853\,
            I => \N__39847\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__39850\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__8455\ : Odrv4
    port map (
            O => \N__39847\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__8454\ : CascadeMux
    port map (
            O => \N__39842\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39833\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39833\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39833\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39827\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__39827\,
            I => \N__39824\
        );

    \I__8448\ : Span4Mux_v
    port map (
            O => \N__39824\,
            I => \N__39820\
        );

    \I__8447\ : InMux
    port map (
            O => \N__39823\,
            I => \N__39817\
        );

    \I__8446\ : Odrv4
    port map (
            O => \N__39820\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39817\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__39812\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39803\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39808\,
            I => \N__39803\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39803\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__8440\ : CascadeMux
    port map (
            O => \N__39800\,
            I => \N__39796\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39793\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39790\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__39793\,
            I => \N__39784\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39790\,
            I => \N__39784\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39789\,
            I => \N__39781\
        );

    \I__8434\ : Span4Mux_v
    port map (
            O => \N__39784\,
            I => \N__39778\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__39781\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8432\ : Odrv4
    port map (
            O => \N__39778\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39768\
        );

    \I__8430\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39765\
        );

    \I__8429\ : CascadeMux
    port map (
            O => \N__39771\,
            I => \N__39761\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39768\,
            I => \N__39758\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__39765\,
            I => \N__39755\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39764\,
            I => \N__39750\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39750\
        );

    \I__8424\ : Span4Mux_v
    port map (
            O => \N__39758\,
            I => \N__39743\
        );

    \I__8423\ : Span4Mux_v
    port map (
            O => \N__39755\,
            I => \N__39743\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39750\,
            I => \N__39743\
        );

    \I__8421\ : Odrv4
    port map (
            O => \N__39743\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39740\,
            I => \N__39736\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39739\,
            I => \N__39733\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39736\,
            I => \N__39727\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__39733\,
            I => \N__39727\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39724\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__39727\,
            I => \N__39721\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39724\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8413\ : Odrv4
    port map (
            O => \N__39721\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39716\,
            I => \N__39712\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39715\,
            I => \N__39707\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__39712\,
            I => \N__39704\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39711\,
            I => \N__39699\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39699\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__39707\,
            I => \N__39696\
        );

    \I__8406\ : Span4Mux_v
    port map (
            O => \N__39704\,
            I => \N__39691\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__39699\,
            I => \N__39691\
        );

    \I__8404\ : Odrv12
    port map (
            O => \N__39696\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8403\ : Odrv4
    port map (
            O => \N__39691\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39686\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__39683\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39674\
        );

    \I__8399\ : InMux
    port map (
            O => \N__39679\,
            I => \N__39674\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__39674\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__8397\ : CascadeMux
    port map (
            O => \N__39671\,
            I => \N__39666\
        );

    \I__8396\ : InMux
    port map (
            O => \N__39670\,
            I => \N__39660\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39669\,
            I => \N__39660\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39655\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39655\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__39660\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__39655\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39650\,
            I => \N__39641\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39641\
        );

    \I__8388\ : InMux
    port map (
            O => \N__39648\,
            I => \N__39641\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39641\,
            I => \N__39638\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__39638\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39635\,
            I => \N__39626\
        );

    \I__8384\ : InMux
    port map (
            O => \N__39634\,
            I => \N__39626\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39626\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__39626\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__8381\ : CascadeMux
    port map (
            O => \N__39623\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39620\,
            I => \N__39617\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__39614\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39607\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39604\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__39607\,
            I => \N__39601\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__39604\,
            I => \N__39598\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__39601\,
            I => \N__39595\
        );

    \I__8372\ : Span4Mux_h
    port map (
            O => \N__39598\,
            I => \N__39588\
        );

    \I__8371\ : Span4Mux_v
    port map (
            O => \N__39595\,
            I => \N__39588\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39594\,
            I => \N__39583\
        );

    \I__8369\ : InMux
    port map (
            O => \N__39593\,
            I => \N__39583\
        );

    \I__8368\ : Span4Mux_v
    port map (
            O => \N__39588\,
            I => \N__39580\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__39583\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8366\ : Odrv4
    port map (
            O => \N__39580\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8365\ : CEMux
    port map (
            O => \N__39575\,
            I => \N__39571\
        );

    \I__8364\ : CEMux
    port map (
            O => \N__39574\,
            I => \N__39566\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__39571\,
            I => \N__39563\
        );

    \I__8362\ : CEMux
    port map (
            O => \N__39570\,
            I => \N__39560\
        );

    \I__8361\ : CEMux
    port map (
            O => \N__39569\,
            I => \N__39557\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39566\,
            I => \N__39554\
        );

    \I__8359\ : Span4Mux_v
    port map (
            O => \N__39563\,
            I => \N__39547\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__39560\,
            I => \N__39547\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__39557\,
            I => \N__39547\
        );

    \I__8356\ : Span4Mux_v
    port map (
            O => \N__39554\,
            I => \N__39542\
        );

    \I__8355\ : Span4Mux_v
    port map (
            O => \N__39547\,
            I => \N__39542\
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__39542\,
            I => \delay_measurement_inst.delay_hc_timer.N_202_i\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39525\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39525\
        );

    \I__8351\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39525\
        );

    \I__8350\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39525\
        );

    \I__8349\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39496\
        );

    \I__8348\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39496\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__39525\,
            I => \N__39493\
        );

    \I__8346\ : InMux
    port map (
            O => \N__39524\,
            I => \N__39484\
        );

    \I__8345\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39484\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39522\,
            I => \N__39484\
        );

    \I__8343\ : InMux
    port map (
            O => \N__39521\,
            I => \N__39484\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39520\,
            I => \N__39475\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39475\
        );

    \I__8340\ : InMux
    port map (
            O => \N__39518\,
            I => \N__39475\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39475\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39466\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39466\
        );

    \I__8336\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39466\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39466\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39457\
        );

    \I__8333\ : InMux
    port map (
            O => \N__39511\,
            I => \N__39457\
        );

    \I__8332\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39457\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39457\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39508\,
            I => \N__39448\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39448\
        );

    \I__8328\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39448\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39448\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39439\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39503\,
            I => \N__39439\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39502\,
            I => \N__39439\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39501\,
            I => \N__39439\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39496\,
            I => \N__39436\
        );

    \I__8321\ : Span4Mux_h
    port map (
            O => \N__39493\,
            I => \N__39431\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__39484\,
            I => \N__39431\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39475\,
            I => \N__39418\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__39466\,
            I => \N__39418\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39457\,
            I => \N__39418\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__39448\,
            I => \N__39418\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__39439\,
            I => \N__39418\
        );

    \I__8314\ : Span4Mux_h
    port map (
            O => \N__39436\,
            I => \N__39418\
        );

    \I__8313\ : Span4Mux_v
    port map (
            O => \N__39431\,
            I => \N__39415\
        );

    \I__8312\ : Span4Mux_v
    port map (
            O => \N__39418\,
            I => \N__39412\
        );

    \I__8311\ : Odrv4
    port map (
            O => \N__39415\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8310\ : Odrv4
    port map (
            O => \N__39412\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8309\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39402\
        );

    \I__8308\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39397\
        );

    \I__8307\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39397\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__39402\,
            I => \N__39391\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__39397\,
            I => \N__39391\
        );

    \I__8304\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39388\
        );

    \I__8303\ : Span12Mux_v
    port map (
            O => \N__39391\,
            I => \N__39385\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__39388\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8301\ : Odrv12
    port map (
            O => \N__39385\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39376\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39379\,
            I => \N__39372\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__39376\,
            I => \N__39369\
        );

    \I__8297\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39366\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39363\
        );

    \I__8295\ : Span4Mux_h
    port map (
            O => \N__39369\,
            I => \N__39360\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__39366\,
            I => \N__39357\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__39363\,
            I => \N__39352\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__39360\,
            I => \N__39352\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__39357\,
            I => \N__39349\
        );

    \I__8290\ : Span4Mux_v
    port map (
            O => \N__39352\,
            I => \N__39346\
        );

    \I__8289\ : Sp12to4
    port map (
            O => \N__39349\,
            I => \N__39343\
        );

    \I__8288\ : Odrv4
    port map (
            O => \N__39346\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8287\ : Odrv12
    port map (
            O => \N__39343\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8286\ : InMux
    port map (
            O => \N__39338\,
            I => \N__39335\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__39335\,
            I => \N__39331\
        );

    \I__8284\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39327\
        );

    \I__8283\ : Span4Mux_v
    port map (
            O => \N__39331\,
            I => \N__39324\
        );

    \I__8282\ : InMux
    port map (
            O => \N__39330\,
            I => \N__39321\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__39327\,
            I => \N__39318\
        );

    \I__8280\ : Span4Mux_v
    port map (
            O => \N__39324\,
            I => \N__39315\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39321\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__39318\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__39315\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8276\ : InMux
    port map (
            O => \N__39308\,
            I => \N__39304\
        );

    \I__8275\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39300\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__39304\,
            I => \N__39297\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39303\,
            I => \N__39294\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__39300\,
            I => \N__39291\
        );

    \I__8271\ : Span12Mux_v
    port map (
            O => \N__39297\,
            I => \N__39288\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__39294\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__39291\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__8268\ : Odrv12
    port map (
            O => \N__39288\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39281\,
            I => \N__39276\
        );

    \I__8266\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39273\
        );

    \I__8265\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39270\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__39276\,
            I => \N__39267\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__39273\,
            I => \N__39264\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__39270\,
            I => \N__39259\
        );

    \I__8261\ : Span4Mux_v
    port map (
            O => \N__39267\,
            I => \N__39259\
        );

    \I__8260\ : Odrv12
    port map (
            O => \N__39264\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__39259\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8258\ : InMux
    port map (
            O => \N__39254\,
            I => \N__39248\
        );

    \I__8257\ : InMux
    port map (
            O => \N__39253\,
            I => \N__39243\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39243\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39240\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__39248\,
            I => \N__39235\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__39243\,
            I => \N__39235\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__39240\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__8251\ : Odrv12
    port map (
            O => \N__39235\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__8250\ : InMux
    port map (
            O => \N__39230\,
            I => \N__39220\
        );

    \I__8249\ : InMux
    port map (
            O => \N__39229\,
            I => \N__39220\
        );

    \I__8248\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39220\
        );

    \I__8247\ : InMux
    port map (
            O => \N__39227\,
            I => \N__39216\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__39220\,
            I => \N__39211\
        );

    \I__8245\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39208\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__39216\,
            I => \N__39205\
        );

    \I__8243\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39202\
        );

    \I__8242\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39199\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__39211\,
            I => \N__39196\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__39208\,
            I => \N__39188\
        );

    \I__8239\ : Span4Mux_h
    port map (
            O => \N__39205\,
            I => \N__39188\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__39202\,
            I => \N__39188\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__39199\,
            I => \N__39183\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__39196\,
            I => \N__39183\
        );

    \I__8235\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39180\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__39188\,
            I => state_3
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__39183\,
            I => state_3
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__39180\,
            I => state_3
        );

    \I__8231\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39169\
        );

    \I__8230\ : InMux
    port map (
            O => \N__39172\,
            I => \N__39163\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__39169\,
            I => \N__39160\
        );

    \I__8228\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39157\
        );

    \I__8227\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39152\
        );

    \I__8226\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39152\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__39163\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__39160\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__39157\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__39152\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__8221\ : IoInMux
    port map (
            O => \N__39143\,
            I => \N__39140\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__39140\,
            I => \N__39137\
        );

    \I__8219\ : Span4Mux_s2_v
    port map (
            O => \N__39137\,
            I => \N__39134\
        );

    \I__8218\ : Span4Mux_v
    port map (
            O => \N__39134\,
            I => \N__39131\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__39131\,
            I => \N__39128\
        );

    \I__8216\ : Span4Mux_v
    port map (
            O => \N__39128\,
            I => \N__39124\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39121\
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__39124\,
            I => \T01_c\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__39121\,
            I => \T01_c\
        );

    \I__8212\ : InMux
    port map (
            O => \N__39116\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__8211\ : InMux
    port map (
            O => \N__39113\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__8210\ : InMux
    port map (
            O => \N__39110\,
            I => \N__39107\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__39107\,
            I => \N__39103\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39099\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__39103\,
            I => \N__39096\
        );

    \I__8206\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39093\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__39099\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__39096\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__39093\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8202\ : InMux
    port map (
            O => \N__39086\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__8201\ : InMux
    port map (
            O => \N__39083\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__39080\,
            I => \N__39076\
        );

    \I__8199\ : CascadeMux
    port map (
            O => \N__39079\,
            I => \N__39072\
        );

    \I__8198\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8197\ : InMux
    port map (
            O => \N__39075\,
            I => \N__39067\
        );

    \I__8196\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39064\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__39067\,
            I => \N__39061\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__39064\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8193\ : Odrv4
    port map (
            O => \N__39061\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8192\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39053\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__39053\,
            I => \N__39050\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__39050\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__8189\ : CascadeMux
    port map (
            O => \N__39047\,
            I => \N__39044\
        );

    \I__8188\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39041\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__39041\,
            I => \N__39038\
        );

    \I__8186\ : Span4Mux_h
    port map (
            O => \N__39038\,
            I => \N__39035\
        );

    \I__8185\ : Span4Mux_v
    port map (
            O => \N__39035\,
            I => \N__39032\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__39032\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__8183\ : InMux
    port map (
            O => \N__39029\,
            I => \N__39026\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__39026\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__8181\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39020\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__39020\,
            I => \N__39017\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__39017\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__8178\ : CascadeMux
    port map (
            O => \N__39014\,
            I => \N__39011\
        );

    \I__8177\ : InMux
    port map (
            O => \N__39011\,
            I => \N__39008\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__39008\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__8175\ : InMux
    port map (
            O => \N__39005\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__8174\ : InMux
    port map (
            O => \N__39002\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38999\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38996\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__8171\ : InMux
    port map (
            O => \N__38993\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38990\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__8169\ : CascadeMux
    port map (
            O => \N__38987\,
            I => \N__38984\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38981\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__38981\,
            I => \N__38977\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38974\
        );

    \I__8165\ : Span4Mux_v
    port map (
            O => \N__38977\,
            I => \N__38968\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38974\,
            I => \N__38968\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38965\
        );

    \I__8162\ : Span4Mux_h
    port map (
            O => \N__38968\,
            I => \N__38962\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38965\,
            I => \N__38959\
        );

    \I__8160\ : Odrv4
    port map (
            O => \N__38962\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8159\ : Odrv12
    port map (
            O => \N__38959\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38954\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__8157\ : InMux
    port map (
            O => \N__38951\,
            I => \bfn_16_11_0_\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38948\,
            I => \N__38945\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__38945\,
            I => \N__38942\
        );

    \I__8154\ : Span4Mux_h
    port map (
            O => \N__38942\,
            I => \N__38937\
        );

    \I__8153\ : InMux
    port map (
            O => \N__38941\,
            I => \N__38932\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38940\,
            I => \N__38932\
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__38937\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__38932\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38927\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38918\
        );

    \I__8146\ : Span4Mux_v
    port map (
            O => \N__38918\,
            I => \N__38915\
        );

    \I__8145\ : Odrv4
    port map (
            O => \N__38915\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__38912\,
            I => \N__38908\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38905\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38908\,
            I => \N__38901\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__38905\,
            I => \N__38898\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38895\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__38901\,
            I => \N__38892\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__38898\,
            I => \N__38889\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38895\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__38892\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__38889\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38882\,
            I => \bfn_16_9_0_\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38879\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38876\,
            I => \N__38873\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38873\,
            I => \N__38868\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38865\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38862\
        );

    \I__8128\ : Odrv4
    port map (
            O => \N__38868\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38865\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__38862\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__8125\ : InMux
    port map (
            O => \N__38855\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__8124\ : InMux
    port map (
            O => \N__38852\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38849\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38846\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38843\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38840\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38837\,
            I => \bfn_16_10_0_\
        );

    \I__8118\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38831\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38831\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38823\
        );

    \I__8115\ : CascadeMux
    port map (
            O => \N__38827\,
            I => \N__38820\
        );

    \I__8114\ : InMux
    port map (
            O => \N__38826\,
            I => \N__38817\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__38823\,
            I => \N__38814\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38820\,
            I => \N__38811\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38817\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8110\ : Odrv4
    port map (
            O => \N__38814\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__38811\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38804\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__8107\ : InMux
    port map (
            O => \N__38801\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38798\,
            I => \N__38795\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__38795\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38792\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38789\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38786\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38780\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38780\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38777\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__8098\ : InMux
    port map (
            O => \N__38774\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38768\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38768\,
            I => \N__38765\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__38765\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__38762\,
            I => \N__38759\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38756\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38756\,
            I => \N__38753\
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__38753\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__38750\,
            I => \N__38747\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38744\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38744\,
            I => \N__38741\
        );

    \I__8087\ : Odrv12
    port map (
            O => \N__38741\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__38738\,
            I => \N__38735\
        );

    \I__8085\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38732\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38732\,
            I => \N__38729\
        );

    \I__8083\ : Odrv12
    port map (
            O => \N__38729\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__38726\,
            I => \N__38723\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38723\,
            I => \N__38720\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__38720\,
            I => \N__38717\
        );

    \I__8079\ : Odrv4
    port map (
            O => \N__38717\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38708\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__38708\,
            I => \N__38705\
        );

    \I__8075\ : Span4Mux_h
    port map (
            O => \N__38705\,
            I => \N__38702\
        );

    \I__8074\ : Odrv4
    port map (
            O => \N__38702\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__38699\,
            I => \N__38696\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38696\,
            I => \N__38693\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38693\,
            I => \N__38690\
        );

    \I__8070\ : Sp12to4
    port map (
            O => \N__38690\,
            I => \N__38687\
        );

    \I__8069\ : Odrv12
    port map (
            O => \N__38687\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__38684\,
            I => \N__38681\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__38678\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__38675\,
            I => \N__38671\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38666\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38666\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38666\,
            I => \N__38662\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38665\,
            I => \N__38659\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__38662\,
            I => \N__38656\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38659\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__38656\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__38651\,
            I => \N__38647\
        );

    \I__8056\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38642\
        );

    \I__8055\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38642\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__38642\,
            I => \N__38638\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38635\
        );

    \I__8052\ : Span4Mux_v
    port map (
            O => \N__38638\,
            I => \N__38632\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__38635\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8050\ : Odrv4
    port map (
            O => \N__38632\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8049\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38621\
        );

    \I__8048\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38621\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__38621\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38615\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__38615\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__8044\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38609\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38609\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__8042\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38603\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__38603\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__8040\ : CascadeMux
    port map (
            O => \N__38600\,
            I => \N__38596\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__38599\,
            I => \N__38593\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38589\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38586\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38583\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__38589\,
            I => \N__38579\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__38586\,
            I => \N__38574\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__38583\,
            I => \N__38574\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38571\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__38579\,
            I => \N__38568\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__38574\,
            I => \N__38565\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__38571\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8028\ : Odrv4
    port map (
            O => \N__38568\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8027\ : Odrv4
    port map (
            O => \N__38565\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8026\ : CascadeMux
    port map (
            O => \N__38558\,
            I => \N__38554\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38550\
        );

    \I__8024\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38547\
        );

    \I__8023\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38544\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38550\,
            I => \N__38538\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38538\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__38544\,
            I => \N__38535\
        );

    \I__8019\ : InMux
    port map (
            O => \N__38543\,
            I => \N__38532\
        );

    \I__8018\ : Span4Mux_v
    port map (
            O => \N__38538\,
            I => \N__38529\
        );

    \I__8017\ : Span4Mux_v
    port map (
            O => \N__38535\,
            I => \N__38526\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38532\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8015\ : Odrv4
    port map (
            O => \N__38529\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8014\ : Odrv4
    port map (
            O => \N__38526\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8013\ : CascadeMux
    port map (
            O => \N__38519\,
            I => \N__38516\
        );

    \I__8012\ : InMux
    port map (
            O => \N__38516\,
            I => \N__38512\
        );

    \I__8011\ : InMux
    port map (
            O => \N__38515\,
            I => \N__38509\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38512\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__38509\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38501\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__38501\,
            I => \N__38498\
        );

    \I__8006\ : Span4Mux_v
    port map (
            O => \N__38498\,
            I => \N__38495\
        );

    \I__8005\ : Odrv4
    port map (
            O => \N__38495\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__8004\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38489\,
            I => \N__38486\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__38486\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__8001\ : InMux
    port map (
            O => \N__38483\,
            I => \N__38480\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__38480\,
            I => \N__38477\
        );

    \I__7999\ : Odrv12
    port map (
            O => \N__38477\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__7998\ : InMux
    port map (
            O => \N__38474\,
            I => \N__38469\
        );

    \I__7997\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38466\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38463\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38469\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__38466\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__38463\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7992\ : CascadeMux
    port map (
            O => \N__38456\,
            I => \N__38452\
        );

    \I__7991\ : CascadeMux
    port map (
            O => \N__38455\,
            I => \N__38448\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38445\
        );

    \I__7989\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38442\
        );

    \I__7988\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38439\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__38445\,
            I => \N__38436\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38442\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__38439\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__38436\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7983\ : CascadeMux
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38423\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__38423\,
            I => \N__38420\
        );

    \I__7980\ : Span4Mux_v
    port map (
            O => \N__38420\,
            I => \N__38417\
        );

    \I__7979\ : Odrv4
    port map (
            O => \N__38417\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__7978\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38411\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__38411\,
            I => \N__38408\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__38408\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38400\
        );

    \I__7974\ : InMux
    port map (
            O => \N__38404\,
            I => \N__38395\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38395\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38400\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__38395\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__7970\ : CascadeMux
    port map (
            O => \N__38390\,
            I => \N__38385\
        );

    \I__7969\ : InMux
    port map (
            O => \N__38389\,
            I => \N__38382\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38377\
        );

    \I__7967\ : InMux
    port map (
            O => \N__38385\,
            I => \N__38377\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__38382\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__38377\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__38372\,
            I => \N__38369\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38369\,
            I => \N__38366\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__38363\,
            I => \N__38360\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__38360\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__7959\ : InMux
    port map (
            O => \N__38357\,
            I => \N__38354\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__38354\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__38351\,
            I => \N__38348\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38345\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__38345\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__7954\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38338\
        );

    \I__7953\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38335\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__38338\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__38335\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__7950\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__38327\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__7948\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38321\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__38321\,
            I => \N__38318\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__38318\,
            I => \N__38315\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__38315\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__38312\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__7943\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38306\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__38306\,
            I => \N__38303\
        );

    \I__7941\ : Odrv12
    port map (
            O => \N__38303\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__7940\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38296\
        );

    \I__7939\ : InMux
    port map (
            O => \N__38299\,
            I => \N__38293\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__38296\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__38293\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__7936\ : InMux
    port map (
            O => \N__38288\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__7935\ : InMux
    port map (
            O => \N__38285\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__7934\ : InMux
    port map (
            O => \N__38282\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__7933\ : InMux
    port map (
            O => \N__38279\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__7932\ : InMux
    port map (
            O => \N__38276\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38273\,
            I => \N__38270\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__38270\,
            I => \N__38267\
        );

    \I__7929\ : Span4Mux_v
    port map (
            O => \N__38267\,
            I => \N__38264\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__38264\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__7927\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38256\
        );

    \I__7926\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38251\
        );

    \I__7925\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38251\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__38256\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__38251\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__38246\,
            I => \N__38243\
        );

    \I__7921\ : InMux
    port map (
            O => \N__38243\,
            I => \N__38236\
        );

    \I__7920\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38236\
        );

    \I__7919\ : InMux
    port map (
            O => \N__38241\,
            I => \N__38233\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__38236\,
            I => \N__38230\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__38233\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__38230\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__38225\,
            I => \N__38222\
        );

    \I__7914\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38219\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__38219\,
            I => \N__38216\
        );

    \I__7912\ : Span4Mux_v
    port map (
            O => \N__38216\,
            I => \N__38213\
        );

    \I__7911\ : Odrv4
    port map (
            O => \N__38213\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__7910\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38204\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38204\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__38204\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__7907\ : CascadeMux
    port map (
            O => \N__38201\,
            I => \N__38198\
        );

    \I__7906\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38192\
        );

    \I__7905\ : InMux
    port map (
            O => \N__38197\,
            I => \N__38192\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__38192\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38189\,
            I => \bfn_15_19_0_\
        );

    \I__7902\ : InMux
    port map (
            O => \N__38186\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38183\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__7900\ : InMux
    port map (
            O => \N__38180\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__7899\ : InMux
    port map (
            O => \N__38177\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__7898\ : InMux
    port map (
            O => \N__38174\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__7897\ : InMux
    port map (
            O => \N__38171\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__7896\ : InMux
    port map (
            O => \N__38168\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38165\,
            I => \bfn_15_20_0_\
        );

    \I__7894\ : InMux
    port map (
            O => \N__38162\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__7893\ : InMux
    port map (
            O => \N__38159\,
            I => \bfn_15_18_0_\
        );

    \I__7892\ : InMux
    port map (
            O => \N__38156\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38153\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__7890\ : InMux
    port map (
            O => \N__38150\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__7889\ : InMux
    port map (
            O => \N__38147\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38144\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__7887\ : InMux
    port map (
            O => \N__38141\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__7886\ : InMux
    port map (
            O => \N__38138\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__7885\ : InMux
    port map (
            O => \N__38135\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__7884\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38108\
        );

    \I__7883\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38108\
        );

    \I__7882\ : InMux
    port map (
            O => \N__38130\,
            I => \N__38108\
        );

    \I__7881\ : InMux
    port map (
            O => \N__38129\,
            I => \N__38108\
        );

    \I__7880\ : InMux
    port map (
            O => \N__38128\,
            I => \N__38099\
        );

    \I__7879\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38099\
        );

    \I__7878\ : InMux
    port map (
            O => \N__38126\,
            I => \N__38099\
        );

    \I__7877\ : InMux
    port map (
            O => \N__38125\,
            I => \N__38099\
        );

    \I__7876\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38076\
        );

    \I__7875\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38076\
        );

    \I__7874\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38076\
        );

    \I__7873\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38076\
        );

    \I__7872\ : InMux
    port map (
            O => \N__38120\,
            I => \N__38067\
        );

    \I__7871\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38067\
        );

    \I__7870\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38067\
        );

    \I__7869\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38067\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__38108\,
            I => \N__38062\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__38099\,
            I => \N__38062\
        );

    \I__7866\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38053\
        );

    \I__7865\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38053\
        );

    \I__7864\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38053\
        );

    \I__7863\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38053\
        );

    \I__7862\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38048\
        );

    \I__7861\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38048\
        );

    \I__7860\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38039\
        );

    \I__7859\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38039\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38039\
        );

    \I__7857\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38039\
        );

    \I__7856\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38030\
        );

    \I__7855\ : InMux
    port map (
            O => \N__38087\,
            I => \N__38030\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38086\,
            I => \N__38030\
        );

    \I__7853\ : InMux
    port map (
            O => \N__38085\,
            I => \N__38030\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__38076\,
            I => \N__38025\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__38067\,
            I => \N__38025\
        );

    \I__7850\ : Span4Mux_v
    port map (
            O => \N__38062\,
            I => \N__38014\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__38053\,
            I => \N__38014\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__38048\,
            I => \N__38014\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__38039\,
            I => \N__38014\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__38030\,
            I => \N__38014\
        );

    \I__7845\ : Span4Mux_v
    port map (
            O => \N__38025\,
            I => \N__38009\
        );

    \I__7844\ : Span4Mux_v
    port map (
            O => \N__38014\,
            I => \N__38009\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__38009\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7842\ : InMux
    port map (
            O => \N__38006\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__7841\ : CEMux
    port map (
            O => \N__38003\,
            I => \N__37998\
        );

    \I__7840\ : CEMux
    port map (
            O => \N__38002\,
            I => \N__37995\
        );

    \I__7839\ : CEMux
    port map (
            O => \N__38001\,
            I => \N__37992\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37998\,
            I => \N__37988\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__37995\,
            I => \N__37983\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37992\,
            I => \N__37983\
        );

    \I__7835\ : CEMux
    port map (
            O => \N__37991\,
            I => \N__37980\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__37988\,
            I => \N__37973\
        );

    \I__7833\ : Span4Mux_v
    port map (
            O => \N__37983\,
            I => \N__37973\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__37980\,
            I => \N__37973\
        );

    \I__7831\ : Span4Mux_v
    port map (
            O => \N__37973\,
            I => \N__37970\
        );

    \I__7830\ : Span4Mux_h
    port map (
            O => \N__37970\,
            I => \N__37967\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__37967\,
            I => \current_shift_inst.timer_s1.N_168_i\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37964\,
            I => \bfn_15_17_0_\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37961\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37958\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__7825\ : InMux
    port map (
            O => \N__37955\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37952\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37949\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__7822\ : InMux
    port map (
            O => \N__37946\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37943\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37940\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37937\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37934\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37931\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37928\,
            I => \bfn_15_16_0_\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37925\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37922\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37919\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37916\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37913\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37910\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37907\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37904\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37901\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37898\,
            I => \bfn_15_15_0_\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37895\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37892\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37889\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37886\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__7801\ : InMux
    port map (
            O => \N__37883\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37880\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37877\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37874\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37871\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37868\,
            I => \bfn_15_14_0_\
        );

    \I__7795\ : InMux
    port map (
            O => \N__37865\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__37862\,
            I => \N__37859\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37856\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__7791\ : Odrv4
    port map (
            O => \N__37853\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37844\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__37844\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37838\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37838\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37832\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37832\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__7783\ : CascadeMux
    port map (
            O => \N__37829\,
            I => \N__37826\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37823\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37823\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__37820\,
            I => \N__37817\
        );

    \I__7779\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37814\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__37814\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__37811\,
            I => \N__37808\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37805\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__37805\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37802\,
            I => \N__37799\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37799\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37796\,
            I => \bfn_15_13_0_\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__37793\,
            I => \N__37790\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37787\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37787\,
            I => \N__37784\
        );

    \I__7768\ : Odrv4
    port map (
            O => \N__37784\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37781\,
            I => \N__37778\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37778\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37775\,
            I => \N__37772\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37772\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37766\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37766\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__37763\,
            I => \N__37760\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37757\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__37757\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37751\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37751\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__37748\,
            I => \N__37745\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37742\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__37742\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__7753\ : CascadeMux
    port map (
            O => \N__37739\,
            I => \N__37736\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37733\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37733\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37727\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__37727\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__37724\,
            I => \N__37721\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37718\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__37718\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__7745\ : CascadeMux
    port map (
            O => \N__37715\,
            I => \N__37712\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37712\,
            I => \N__37709\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__37709\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__7742\ : CascadeMux
    port map (
            O => \N__37706\,
            I => \N__37703\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37700\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__37700\,
            I => \N__37697\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__37697\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__37694\,
            I => \N__37691\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37688\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37688\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__37685\,
            I => \N__37682\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37679\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__37679\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37676\,
            I => \N__37673\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__37673\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__37670\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__7729\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37661\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37666\,
            I => \N__37658\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37665\,
            I => \N__37653\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37653\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37661\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__37658\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__37653\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__7722\ : CascadeMux
    port map (
            O => \N__37646\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__37643\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__7720\ : CascadeMux
    port map (
            O => \N__37640\,
            I => \N__37637\
        );

    \I__7719\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37633\
        );

    \I__7718\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37630\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37627\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__37630\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__7715\ : Odrv4
    port map (
            O => \N__37627\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__7714\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37619\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__37619\,
            I => \N__37616\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__37616\,
            I => \N__37612\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37615\,
            I => \N__37609\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__37612\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__37609\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7708\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37601\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__37601\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__37598\,
            I => \N__37595\
        );

    \I__7705\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37592\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37587\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__37591\,
            I => \N__37584\
        );

    \I__7702\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37580\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__37587\,
            I => \N__37577\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37574\
        );

    \I__7699\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37571\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__37580\,
            I => \N__37568\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__37577\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__37574\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__37571\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__7694\ : Odrv12
    port map (
            O => \N__37568\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__7693\ : CascadeMux
    port map (
            O => \N__37559\,
            I => \N__37556\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37553\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37553\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37550\,
            I => \N__37547\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__37547\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__7688\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37538\
        );

    \I__7686\ : Span4Mux_v
    port map (
            O => \N__37538\,
            I => \N__37535\
        );

    \I__7685\ : Odrv4
    port map (
            O => \N__37535\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__37532\,
            I => \N__37529\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37529\,
            I => \N__37526\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__37526\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__37520\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__7679\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__37514\,
            I => \N__37511\
        );

    \I__7677\ : Odrv4
    port map (
            O => \N__37511\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__7676\ : CascadeMux
    port map (
            O => \N__37508\,
            I => \N__37505\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37505\,
            I => \N__37502\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37502\,
            I => \N__37499\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__37499\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37490\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__37490\,
            I => \N__37487\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__37487\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__7668\ : CascadeMux
    port map (
            O => \N__37484\,
            I => \N__37481\
        );

    \I__7667\ : InMux
    port map (
            O => \N__37481\,
            I => \N__37478\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__7665\ : Span4Mux_h
    port map (
            O => \N__37475\,
            I => \N__37472\
        );

    \I__7664\ : Odrv4
    port map (
            O => \N__37472\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__7663\ : CascadeMux
    port map (
            O => \N__37469\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7661\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__37460\,
            I => \N__37457\
        );

    \I__7659\ : Odrv12
    port map (
            O => \N__37457\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__37454\,
            I => \N__37451\
        );

    \I__7657\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37448\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__37448\,
            I => \N__37445\
        );

    \I__7655\ : Span4Mux_h
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7654\ : Span4Mux_v
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__37439\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\
        );

    \I__7652\ : IoInMux
    port map (
            O => \N__37436\,
            I => \N__37410\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37435\,
            I => \N__37393\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37393\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37393\
        );

    \I__7648\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37393\
        );

    \I__7647\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37384\
        );

    \I__7646\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37384\
        );

    \I__7645\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37384\
        );

    \I__7644\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37384\
        );

    \I__7643\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37377\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37377\
        );

    \I__7641\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37377\
        );

    \I__7640\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37368\
        );

    \I__7639\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37368\
        );

    \I__7638\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37368\
        );

    \I__7637\ : InMux
    port map (
            O => \N__37421\,
            I => \N__37368\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37420\,
            I => \N__37359\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37359\
        );

    \I__7634\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37359\
        );

    \I__7633\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37359\
        );

    \I__7632\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37350\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37415\,
            I => \N__37350\
        );

    \I__7630\ : InMux
    port map (
            O => \N__37414\,
            I => \N__37350\
        );

    \I__7629\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37350\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__37410\,
            I => \N__37347\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37344\
        );

    \I__7626\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37337\
        );

    \I__7625\ : InMux
    port map (
            O => \N__37407\,
            I => \N__37337\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37406\,
            I => \N__37337\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37328\
        );

    \I__7622\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37328\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37328\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37402\,
            I => \N__37328\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__37393\,
            I => \N__37323\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__37384\,
            I => \N__37323\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37314\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37368\,
            I => \N__37314\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37359\,
            I => \N__37314\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__37350\,
            I => \N__37314\
        );

    \I__7613\ : Span4Mux_s1_v
    port map (
            O => \N__37347\,
            I => \N__37311\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__37344\,
            I => \N__37308\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37299\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37328\,
            I => \N__37299\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__37323\,
            I => \N__37299\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__37314\,
            I => \N__37299\
        );

    \I__7607\ : Span4Mux_h
    port map (
            O => \N__37311\,
            I => \N__37296\
        );

    \I__7606\ : Span4Mux_v
    port map (
            O => \N__37308\,
            I => \N__37289\
        );

    \I__7605\ : Span4Mux_v
    port map (
            O => \N__37299\,
            I => \N__37289\
        );

    \I__7604\ : Span4Mux_v
    port map (
            O => \N__37296\,
            I => \N__37289\
        );

    \I__7603\ : Odrv4
    port map (
            O => \N__37289\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37280\
        );

    \I__7601\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37280\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__37280\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__37277\,
            I => \N__37274\
        );

    \I__7598\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37270\
        );

    \I__7597\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37264\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__37270\,
            I => \N__37261\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37254\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37268\,
            I => \N__37254\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37267\,
            I => \N__37254\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__37264\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7591\ : Odrv4
    port map (
            O => \N__37261\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__37254\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37244\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__37244\,
            I => \N__37239\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37243\,
            I => \N__37236\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__37242\,
            I => \N__37233\
        );

    \I__7585\ : Span4Mux_v
    port map (
            O => \N__37239\,
            I => \N__37228\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37236\,
            I => \N__37228\
        );

    \I__7583\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37225\
        );

    \I__7582\ : Span4Mux_v
    port map (
            O => \N__37228\,
            I => \N__37222\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__37225\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__37222\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7579\ : CascadeMux
    port map (
            O => \N__37217\,
            I => \N__37214\
        );

    \I__7578\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__37211\,
            I => \N__37208\
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__37208\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__7575\ : CascadeMux
    port map (
            O => \N__37205\,
            I => \N__37202\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37199\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__37199\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__37196\,
            I => \N__37193\
        );

    \I__7571\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37190\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__37181\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__7566\ : CascadeMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__7565\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37172\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__7563\ : Odrv4
    port map (
            O => \N__37169\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__37163\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__7560\ : InMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__7557\ : Odrv4
    port map (
            O => \N__37151\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__7555\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__37136\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__37124\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__7546\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37115\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__37115\,
            I => \N__37112\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__37112\,
            I => \N__37109\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__37109\,
            I => \N__37106\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__37106\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__7541\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37097\
        );

    \I__7539\ : Odrv12
    port map (
            O => \N__37097\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7537\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__7535\ : Odrv12
    port map (
            O => \N__37085\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__7534\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37079\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__37079\,
            I => \N__37076\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__37076\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37073\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28\
        );

    \I__7530\ : InMux
    port map (
            O => \N__37070\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__7529\ : InMux
    port map (
            O => \N__37067\,
            I => \N__37063\
        );

    \I__7528\ : InMux
    port map (
            O => \N__37066\,
            I => \N__37060\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__37063\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__37060\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7525\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37052\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__37052\,
            I => \N__37045\
        );

    \I__7523\ : InMux
    port map (
            O => \N__37051\,
            I => \N__37042\
        );

    \I__7522\ : InMux
    port map (
            O => \N__37050\,
            I => \N__37039\
        );

    \I__7521\ : InMux
    port map (
            O => \N__37049\,
            I => \N__37036\
        );

    \I__7520\ : InMux
    port map (
            O => \N__37048\,
            I => \N__37033\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__37045\,
            I => \N__37030\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__37042\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__37039\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__37036\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__37033\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__37030\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__37019\,
            I => \N__37016\
        );

    \I__7512\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__37013\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df30\
        );

    \I__7510\ : InMux
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__37007\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__7508\ : InMux
    port map (
            O => \N__37004\,
            I => \N__37000\
        );

    \I__7507\ : InMux
    port map (
            O => \N__37003\,
            I => \N__36997\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__37000\,
            I => \N__36994\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__36997\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7504\ : Odrv12
    port map (
            O => \N__36994\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36986\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__36980\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__7499\ : CascadeMux
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7498\ : InMux
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36971\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36965\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__36965\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36962\,
            I => \N__36958\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36955\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36958\,
            I => \N__36952\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__36955\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7490\ : Odrv12
    port map (
            O => \N__36952\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7489\ : CascadeMux
    port map (
            O => \N__36947\,
            I => \N__36944\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36944\,
            I => \N__36941\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36941\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__36938\,
            I => \N__36935\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36932\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36932\,
            I => \N__36929\
        );

    \I__7483\ : Odrv12
    port map (
            O => \N__36929\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36926\,
            I => \N__36922\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36925\,
            I => \N__36919\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__36922\,
            I => \N__36916\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__36919\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7478\ : Odrv12
    port map (
            O => \N__36916\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36908\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36908\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36899\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__36899\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36893\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36893\,
            I => \N__36889\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36886\
        );

    \I__7469\ : Span4Mux_v
    port map (
            O => \N__36889\,
            I => \N__36883\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__36886\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__36883\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36875\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__36875\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36869\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36869\,
            I => \N__36866\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__36866\,
            I => \N__36863\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__36863\,
            I => \N__36860\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__36860\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36857\,
            I => \N__36853\
        );

    \I__7458\ : InMux
    port map (
            O => \N__36856\,
            I => \N__36850\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__36853\,
            I => \N__36847\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36850\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7455\ : Odrv12
    port map (
            O => \N__36847\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__36842\,
            I => \N__36839\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36839\,
            I => \N__36836\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__36836\,
            I => \N__36833\
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__36833\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36826\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36823\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36826\,
            I => \N__36820\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__36823\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7446\ : Odrv12
    port map (
            O => \N__36820\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36812\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36812\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36809\,
            I => \N__36806\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__36806\,
            I => \N__36802\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36805\,
            I => \N__36799\
        );

    \I__7440\ : Span4Mux_v
    port map (
            O => \N__36802\,
            I => \N__36796\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36799\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__36796\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36791\,
            I => \N__36788\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36788\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36782\,
            I => \N__36778\
        );

    \I__7433\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36775\
        );

    \I__7432\ : Span4Mux_v
    port map (
            O => \N__36778\,
            I => \N__36772\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__36775\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__36772\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36761\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36751\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36754\,
            I => \N__36748\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__36751\,
            I => \N__36745\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__36748\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7421\ : Odrv4
    port map (
            O => \N__36745\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7420\ : CascadeMux
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36734\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__36734\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36727\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36730\,
            I => \N__36724\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__36727\,
            I => \N__36721\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__36724\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7413\ : Odrv12
    port map (
            O => \N__36721\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__36716\,
            I => \N__36713\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36710\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__36704\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36697\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36694\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__36697\,
            I => \N__36691\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__36694\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7403\ : Odrv12
    port map (
            O => \N__36691\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__36686\,
            I => \N__36683\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36683\,
            I => \N__36680\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__36680\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36674\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__36674\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36671\,
            I => \N__36667\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36664\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__36667\,
            I => \N__36661\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__36664\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7393\ : Odrv12
    port map (
            O => \N__36661\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7392\ : CascadeMux
    port map (
            O => \N__36656\,
            I => \N__36653\
        );

    \I__7391\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36650\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36650\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__7389\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__36644\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36641\,
            I => \N__36637\
        );

    \I__7386\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36634\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__36637\,
            I => \N__36631\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__36634\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7383\ : Odrv12
    port map (
            O => \N__36631\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7382\ : CascadeMux
    port map (
            O => \N__36626\,
            I => \N__36623\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36620\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__36620\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__7379\ : InMux
    port map (
            O => \N__36617\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36614\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__7377\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36605\
        );

    \I__7376\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36605\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36602\
        );

    \I__7374\ : Odrv12
    port map (
            O => \N__36602\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__7373\ : InMux
    port map (
            O => \N__36599\,
            I => \N__36594\
        );

    \I__7372\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36589\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36589\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__36594\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__36589\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7368\ : CascadeMux
    port map (
            O => \N__36584\,
            I => \N__36581\
        );

    \I__7367\ : InMux
    port map (
            O => \N__36581\,
            I => \N__36574\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36574\
        );

    \I__7365\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36571\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__36574\,
            I => \N__36568\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__36571\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7362\ : Odrv4
    port map (
            O => \N__36568\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__7360\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36554\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36554\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__36554\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__7357\ : CascadeMux
    port map (
            O => \N__36551\,
            I => \N__36548\
        );

    \I__7356\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__36545\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__7354\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36539\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__36539\,
            I => \N__36535\
        );

    \I__7352\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36532\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__36535\,
            I => \N__36529\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36532\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7349\ : Odrv4
    port map (
            O => \N__36529\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__36524\,
            I => \N__36521\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36521\,
            I => \N__36518\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36515\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__36515\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__7344\ : CascadeMux
    port map (
            O => \N__36512\,
            I => \N__36507\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36511\,
            I => \N__36504\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36510\,
            I => \N__36499\
        );

    \I__7341\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36499\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36504\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__36499\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36494\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__36491\,
            I => \N__36486\
        );

    \I__7336\ : InMux
    port map (
            O => \N__36490\,
            I => \N__36483\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36478\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36478\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36483\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__36478\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36473\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__36470\,
            I => \N__36465\
        );

    \I__7329\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36462\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36468\,
            I => \N__36457\
        );

    \I__7327\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36457\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__36462\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__36457\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__7324\ : InMux
    port map (
            O => \N__36452\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__7323\ : InMux
    port map (
            O => \N__36449\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__7322\ : InMux
    port map (
            O => \N__36446\,
            I => \bfn_14_22_0_\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36443\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36440\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__7319\ : InMux
    port map (
            O => \N__36437\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__7318\ : InMux
    port map (
            O => \N__36434\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__7317\ : InMux
    port map (
            O => \N__36431\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__7316\ : InMux
    port map (
            O => \N__36428\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__7315\ : InMux
    port map (
            O => \N__36425\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36422\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__7313\ : InMux
    port map (
            O => \N__36419\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__7312\ : InMux
    port map (
            O => \N__36416\,
            I => \bfn_14_21_0_\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36413\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36410\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__7309\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36402\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36397\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36397\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__36402\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__36397\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7304\ : InMux
    port map (
            O => \N__36392\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__7303\ : InMux
    port map (
            O => \N__36389\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__7302\ : InMux
    port map (
            O => \N__36386\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36383\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__7300\ : InMux
    port map (
            O => \N__36380\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__7299\ : InMux
    port map (
            O => \N__36377\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36374\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36371\,
            I => \bfn_14_20_0_\
        );

    \I__7296\ : InMux
    port map (
            O => \N__36368\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__7295\ : InMux
    port map (
            O => \N__36365\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__7294\ : IoInMux
    port map (
            O => \N__36362\,
            I => \N__36359\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36356\
        );

    \I__7292\ : IoSpan4Mux
    port map (
            O => \N__36356\,
            I => \N__36353\
        );

    \I__7291\ : Span4Mux_s3_v
    port map (
            O => \N__36353\,
            I => \N__36350\
        );

    \I__7290\ : Sp12to4
    port map (
            O => \N__36350\,
            I => \N__36347\
        );

    \I__7289\ : Span12Mux_v
    port map (
            O => \N__36347\,
            I => \N__36344\
        );

    \I__7288\ : Odrv12
    port map (
            O => \N__36344\,
            I => \pll_inst.red_c_i\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__36341\,
            I => \N__36338\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36338\,
            I => \N__36333\
        );

    \I__7285\ : InMux
    port map (
            O => \N__36337\,
            I => \N__36330\
        );

    \I__7284\ : InMux
    port map (
            O => \N__36336\,
            I => \N__36327\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__36333\,
            I => \N__36324\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__36330\,
            I => \N__36321\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__36327\,
            I => \N__36314\
        );

    \I__7280\ : Span12Mux_h
    port map (
            O => \N__36324\,
            I => \N__36314\
        );

    \I__7279\ : Sp12to4
    port map (
            O => \N__36321\,
            I => \N__36314\
        );

    \I__7278\ : Span12Mux_v
    port map (
            O => \N__36314\,
            I => \N__36311\
        );

    \I__7277\ : Odrv12
    port map (
            O => \N__36311\,
            I => \il_max_comp1_D2\
        );

    \I__7276\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__36305\,
            I => \N__36301\
        );

    \I__7274\ : InMux
    port map (
            O => \N__36304\,
            I => \N__36297\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__36301\,
            I => \N__36294\
        );

    \I__7272\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36291\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__36297\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__7270\ : Odrv4
    port map (
            O => \N__36294\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36291\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__7268\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36281\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__36281\,
            I => \N__36277\
        );

    \I__7266\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36273\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__36277\,
            I => \N__36270\
        );

    \I__7264\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36267\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__36273\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7262\ : Odrv4
    port map (
            O => \N__36270\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__36267\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__7260\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36256\
        );

    \I__7259\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36252\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36249\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36246\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__36252\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__7255\ : Odrv4
    port map (
            O => \N__36249\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__36246\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__7253\ : InMux
    port map (
            O => \N__36239\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__7252\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36233\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36233\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7250\ : InMux
    port map (
            O => \N__36230\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__7249\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36224\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__36224\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__7247\ : InMux
    port map (
            O => \N__36221\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__7246\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36215\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__36215\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__7244\ : InMux
    port map (
            O => \N__36212\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__7243\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36206\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__36206\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__7241\ : InMux
    port map (
            O => \N__36203\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__7240\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36197\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__36197\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__7238\ : InMux
    port map (
            O => \N__36194\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36188\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36185\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__36185\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36182\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__36179\,
            I => \N__36176\
        );

    \I__7232\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36173\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__36173\,
            I => \N__36170\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__36170\,
            I => \N__36167\
        );

    \I__7229\ : Odrv4
    port map (
            O => \N__36167\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__7228\ : InMux
    port map (
            O => \N__36164\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__7227\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36158\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__36158\,
            I => \N__36155\
        );

    \I__7225\ : Odrv4
    port map (
            O => \N__36155\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__7224\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__36149\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__7222\ : InMux
    port map (
            O => \N__36146\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__7221\ : InMux
    port map (
            O => \N__36143\,
            I => \N__36140\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36140\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__7219\ : InMux
    port map (
            O => \N__36137\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__7218\ : InMux
    port map (
            O => \N__36134\,
            I => \N__36131\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__36131\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__7216\ : InMux
    port map (
            O => \N__36128\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__7215\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36122\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__36122\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7213\ : InMux
    port map (
            O => \N__36119\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__7212\ : InMux
    port map (
            O => \N__36116\,
            I => \N__36113\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__36113\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7210\ : InMux
    port map (
            O => \N__36110\,
            I => \bfn_14_12_0_\
        );

    \I__7209\ : InMux
    port map (
            O => \N__36107\,
            I => \N__36104\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36104\,
            I => \N__36101\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__36101\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__7206\ : InMux
    port map (
            O => \N__36098\,
            I => \N__36095\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__36095\,
            I => \N__36092\
        );

    \I__7204\ : Span4Mux_v
    port map (
            O => \N__36092\,
            I => \N__36089\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__36089\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__7202\ : InMux
    port map (
            O => \N__36086\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__7201\ : InMux
    port map (
            O => \N__36083\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__7200\ : InMux
    port map (
            O => \N__36080\,
            I => \N__36077\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36074\
        );

    \I__7198\ : Span4Mux_h
    port map (
            O => \N__36074\,
            I => \N__36071\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__36071\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__36068\,
            I => \N__36065\
        );

    \I__7195\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36062\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__36062\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__7193\ : CascadeMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7192\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36053\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__36053\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__7190\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36047\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__36047\,
            I => \N__36044\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__36044\,
            I => \N__36041\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__36041\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__7186\ : InMux
    port map (
            O => \N__36038\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__7185\ : InMux
    port map (
            O => \N__36035\,
            I => \N__36032\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__36032\,
            I => \N__36029\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__36029\,
            I => \N__36026\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__36026\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__7181\ : InMux
    port map (
            O => \N__36023\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__36020\,
            I => \N__36017\
        );

    \I__7179\ : InMux
    port map (
            O => \N__36017\,
            I => \N__36014\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__36014\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__7177\ : InMux
    port map (
            O => \N__36011\,
            I => \N__36008\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__36008\,
            I => \N__36005\
        );

    \I__7175\ : Span4Mux_v
    port map (
            O => \N__36005\,
            I => \N__36002\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__36002\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35999\,
            I => \bfn_14_8_0_\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35993\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__35993\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__7170\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35987\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__35987\,
            I => \N__35984\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__35984\,
            I => \N__35981\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__35981\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35978\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__7165\ : CascadeMux
    port map (
            O => \N__35975\,
            I => \N__35972\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35969\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__35969\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35963\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__35960\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35957\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35954\,
            I => \N__35951\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35951\,
            I => \N__35948\
        );

    \I__7156\ : Odrv4
    port map (
            O => \N__35948\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35945\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35939\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__35939\,
            I => \N__35936\
        );

    \I__7152\ : Odrv4
    port map (
            O => \N__35936\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35933\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__7150\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35927\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__35927\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35924\,
            I => \N__35921\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__35921\,
            I => \N__35918\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__35918\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35915\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35909\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__35909\,
            I => \N__35906\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__35906\,
            I => \N__35903\
        );

    \I__7141\ : Odrv4
    port map (
            O => \N__35903\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35900\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35894\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__35891\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35888\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35882\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__35882\,
            I => \N__35877\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35874\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35868\
        );

    \I__7131\ : Span12Mux_h
    port map (
            O => \N__35877\,
            I => \N__35865\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35874\,
            I => \N__35862\
        );

    \I__7129\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35859\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35856\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35853\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__35868\,
            I => \N__35850\
        );

    \I__7125\ : Odrv12
    port map (
            O => \N__35865\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__35862\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35859\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35856\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35853\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__35850\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7119\ : IoInMux
    port map (
            O => \N__35837\,
            I => \N__35834\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35831\
        );

    \I__7117\ : Odrv12
    port map (
            O => \N__35831\,
            I => s2_phy_c
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__35828\,
            I => \N__35825\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35821\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35818\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35821\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35818\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35808\
        );

    \I__7110\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35805\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35801\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__35808\,
            I => \N__35796\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__35805\,
            I => \N__35796\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__35804\,
            I => \N__35793\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__35801\,
            I => \N__35788\
        );

    \I__7104\ : Span4Mux_v
    port map (
            O => \N__35796\,
            I => \N__35788\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35785\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__35788\,
            I => \N__35782\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35785\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7100\ : Odrv4
    port map (
            O => \N__35782\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7099\ : ClkMux
    port map (
            O => \N__35777\,
            I => \N__35774\
        );

    \I__7098\ : GlobalMux
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__7097\ : gio2CtrlBuf
    port map (
            O => \N__35771\,
            I => delay_hc_input_c_g
        );

    \I__7096\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35765\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35760\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35757\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35754\
        );

    \I__7092\ : Span12Mux_v
    port map (
            O => \N__35760\,
            I => \N__35749\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35757\,
            I => \N__35749\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__35754\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__35749\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__35744\,
            I => \N__35740\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35736\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35740\,
            I => \N__35731\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35731\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__35736\,
            I => \N__35728\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35731\,
            I => \N__35725\
        );

    \I__7082\ : Span12Mux_h
    port map (
            O => \N__35728\,
            I => \N__35721\
        );

    \I__7081\ : Span12Mux_h
    port map (
            O => \N__35725\,
            I => \N__35718\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35715\
        );

    \I__7079\ : Span12Mux_v
    port map (
            O => \N__35721\,
            I => \N__35712\
        );

    \I__7078\ : Span12Mux_v
    port map (
            O => \N__35718\,
            I => \N__35709\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__35715\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__7076\ : Odrv12
    port map (
            O => \N__35712\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__7075\ : Odrv12
    port map (
            O => \N__35709\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35696\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35689\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35689\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35689\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35696\,
            I => \N__35686\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__35689\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7068\ : Odrv12
    port map (
            O => \N__35686\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7067\ : CascadeMux
    port map (
            O => \N__35681\,
            I => \N__35676\
        );

    \I__7066\ : InMux
    port map (
            O => \N__35680\,
            I => \N__35672\
        );

    \I__7065\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35669\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35664\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35664\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__35672\,
            I => \N__35661\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__35669\,
            I => \N__35658\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__35664\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7059\ : Odrv12
    port map (
            O => \N__35661\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__35658\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7057\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35647\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35650\,
            I => \N__35642\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__35647\,
            I => \N__35639\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35636\
        );

    \I__7053\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35633\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35628\
        );

    \I__7051\ : Span12Mux_v
    port map (
            O => \N__35639\,
            I => \N__35628\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__35636\,
            I => \N__35625\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__35633\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7048\ : Odrv12
    port map (
            O => \N__35628\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__35625\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7046\ : IoInMux
    port map (
            O => \N__35618\,
            I => \N__35615\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__7044\ : Span4Mux_s1_v
    port map (
            O => \N__35612\,
            I => \N__35609\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__35609\,
            I => \N__35604\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35599\
        );

    \I__7041\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35599\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__35604\,
            I => s1_phy_c
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__35599\,
            I => s1_phy_c
        );

    \I__7038\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__35591\,
            I => \N__35588\
        );

    \I__7036\ : Odrv12
    port map (
            O => \N__35588\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__7035\ : CascadeMux
    port map (
            O => \N__35585\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__7034\ : IoInMux
    port map (
            O => \N__35582\,
            I => \N__35579\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35579\,
            I => \N__35576\
        );

    \I__7032\ : Odrv12
    port map (
            O => \N__35576\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__7031\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35570\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35565\
        );

    \I__7029\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35562\
        );

    \I__7028\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35559\
        );

    \I__7027\ : Span4Mux_v
    port map (
            O => \N__35565\,
            I => \N__35554\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__35562\,
            I => \N__35554\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35559\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__7024\ : Odrv4
    port map (
            O => \N__35554\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35543\
        );

    \I__7022\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35543\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__35543\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35534\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35534\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35534\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__7017\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35525\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35525\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35525\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__7014\ : CascadeMux
    port map (
            O => \N__35522\,
            I => \N__35519\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35513\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35513\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35513\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__7010\ : IoInMux
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__35507\,
            I => \N__35504\
        );

    \I__7008\ : Span4Mux_s2_v
    port map (
            O => \N__35504\,
            I => \N__35501\
        );

    \I__7007\ : Span4Mux_h
    port map (
            O => \N__35501\,
            I => \N__35498\
        );

    \I__7006\ : Span4Mux_v
    port map (
            O => \N__35498\,
            I => \N__35495\
        );

    \I__7005\ : Span4Mux_v
    port map (
            O => \N__35495\,
            I => \N__35491\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35488\
        );

    \I__7003\ : Odrv4
    port map (
            O => \N__35491\,
            I => \T12_c\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__35488\,
            I => \T12_c\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__35483\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__35477\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__35474\,
            I => \N__35468\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__35473\,
            I => \N__35465\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35462\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35458\
        );

    \I__6994\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35453\
        );

    \I__6993\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35453\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35462\,
            I => \N__35450\
        );

    \I__6991\ : InMux
    port map (
            O => \N__35461\,
            I => \N__35447\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35444\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__35453\,
            I => \N__35441\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__35450\,
            I => \N__35438\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35435\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__35444\,
            I => \N__35432\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__35441\,
            I => \N__35427\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__35438\,
            I => \N__35427\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__35435\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__35432\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__6981\ : Odrv4
    port map (
            O => \N__35427\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__6980\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35417\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__35417\,
            I => \N__35414\
        );

    \I__6978\ : Span4Mux_h
    port map (
            O => \N__35414\,
            I => \N__35411\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__35411\,
            I => \N__35408\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__35408\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__35405\,
            I => \N__35392\
        );

    \I__6974\ : CascadeMux
    port map (
            O => \N__35404\,
            I => \N__35388\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__35403\,
            I => \N__35385\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35377\
        );

    \I__6971\ : CascadeMux
    port map (
            O => \N__35401\,
            I => \N__35372\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__35400\,
            I => \N__35369\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__35399\,
            I => \N__35365\
        );

    \I__6968\ : CascadeMux
    port map (
            O => \N__35398\,
            I => \N__35362\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__35397\,
            I => \N__35359\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__35396\,
            I => \N__35355\
        );

    \I__6965\ : CascadeMux
    port map (
            O => \N__35395\,
            I => \N__35351\
        );

    \I__6964\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35348\
        );

    \I__6963\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35343\
        );

    \I__6962\ : InMux
    port map (
            O => \N__35388\,
            I => \N__35343\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35340\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__35384\,
            I => \N__35327\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__35383\,
            I => \N__35324\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__35382\,
            I => \N__35321\
        );

    \I__6957\ : CascadeMux
    port map (
            O => \N__35381\,
            I => \N__35317\
        );

    \I__6956\ : CascadeMux
    port map (
            O => \N__35380\,
            I => \N__35314\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35311\
        );

    \I__6954\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35302\
        );

    \I__6953\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35302\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35302\
        );

    \I__6951\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35302\
        );

    \I__6950\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35293\
        );

    \I__6949\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35293\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35362\,
            I => \N__35293\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35359\,
            I => \N__35293\
        );

    \I__6946\ : InMux
    port map (
            O => \N__35358\,
            I => \N__35289\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35355\,
            I => \N__35282\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35354\,
            I => \N__35282\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35282\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__35348\,
            I => \N__35279\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__35343\,
            I => \N__35274\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__35340\,
            I => \N__35274\
        );

    \I__6939\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35261\
        );

    \I__6938\ : InMux
    port map (
            O => \N__35338\,
            I => \N__35261\
        );

    \I__6937\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35261\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35261\
        );

    \I__6935\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35261\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35334\,
            I => \N__35261\
        );

    \I__6933\ : InMux
    port map (
            O => \N__35333\,
            I => \N__35254\
        );

    \I__6932\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35254\
        );

    \I__6931\ : InMux
    port map (
            O => \N__35331\,
            I => \N__35254\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35240\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35240\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35240\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35240\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35320\,
            I => \N__35240\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35240\
        );

    \I__6924\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35228\
        );

    \I__6923\ : Span4Mux_v
    port map (
            O => \N__35311\,
            I => \N__35221\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__35302\,
            I => \N__35221\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__35293\,
            I => \N__35221\
        );

    \I__6920\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35218\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__35289\,
            I => \N__35204\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35204\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__35279\,
            I => \N__35204\
        );

    \I__6916\ : Span4Mux_v
    port map (
            O => \N__35274\,
            I => \N__35204\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35204\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35204\
        );

    \I__6913\ : InMux
    port map (
            O => \N__35253\,
            I => \N__35201\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__35240\,
            I => \N__35198\
        );

    \I__6911\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35195\
        );

    \I__6910\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35178\
        );

    \I__6909\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35178\
        );

    \I__6908\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35178\
        );

    \I__6907\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35178\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35178\
        );

    \I__6905\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35178\
        );

    \I__6904\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35178\
        );

    \I__6903\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35178\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35171\
        );

    \I__6901\ : Span4Mux_v
    port map (
            O => \N__35221\,
            I => \N__35166\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__35218\,
            I => \N__35166\
        );

    \I__6899\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35163\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__35204\,
            I => \N__35160\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35151\
        );

    \I__6896\ : Span4Mux_h
    port map (
            O => \N__35198\,
            I => \N__35151\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__35195\,
            I => \N__35151\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__35178\,
            I => \N__35151\
        );

    \I__6893\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35142\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35142\
        );

    \I__6891\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35142\
        );

    \I__6890\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35142\
        );

    \I__6889\ : Odrv12
    port map (
            O => \N__35171\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6888\ : Odrv4
    port map (
            O => \N__35166\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__35163\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__35160\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6885\ : Odrv4
    port map (
            O => \N__35151\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__35142\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6883\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35125\
        );

    \I__6882\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35122\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35116\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__35122\,
            I => \N__35116\
        );

    \I__6879\ : InMux
    port map (
            O => \N__35121\,
            I => \N__35113\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__35116\,
            I => \N__35110\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__35113\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__35110\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__6875\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35102\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__35102\,
            I => \phase_controller_inst1.N_55\
        );

    \I__6873\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35093\
        );

    \I__6872\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35093\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__35093\,
            I => \N__35089\
        );

    \I__6870\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35085\
        );

    \I__6869\ : Span4Mux_h
    port map (
            O => \N__35089\,
            I => \N__35082\
        );

    \I__6868\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35079\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__35085\,
            I => \N__35076\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__35082\,
            I => \N__35073\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__35079\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6864\ : Odrv12
    port map (
            O => \N__35076\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__35073\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6862\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35062\
        );

    \I__6861\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35059\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__35053\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__35059\,
            I => \N__35053\
        );

    \I__6858\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35050\
        );

    \I__6857\ : Span4Mux_s3_v
    port map (
            O => \N__35053\,
            I => \N__35047\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35044\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__35047\,
            I => \N__35041\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__35044\,
            I => \N__35038\
        );

    \I__6853\ : Sp12to4
    port map (
            O => \N__35041\,
            I => \N__35034\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__35038\,
            I => \N__35031\
        );

    \I__6851\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35028\
        );

    \I__6850\ : Span12Mux_v
    port map (
            O => \N__35034\,
            I => \N__35025\
        );

    \I__6849\ : Sp12to4
    port map (
            O => \N__35031\,
            I => \N__35022\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__35028\,
            I => \N__35019\
        );

    \I__6847\ : Span12Mux_v
    port map (
            O => \N__35025\,
            I => \N__35016\
        );

    \I__6846\ : Span12Mux_s7_h
    port map (
            O => \N__35022\,
            I => \N__35011\
        );

    \I__6845\ : Span12Mux_h
    port map (
            O => \N__35019\,
            I => \N__35011\
        );

    \I__6844\ : Span12Mux_h
    port map (
            O => \N__35016\,
            I => \N__35006\
        );

    \I__6843\ : Span12Mux_v
    port map (
            O => \N__35011\,
            I => \N__35006\
        );

    \I__6842\ : Odrv12
    port map (
            O => \N__35006\,
            I => start_stop_c
        );

    \I__6841\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34999\
        );

    \I__6840\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34996\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34993\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34990\
        );

    \I__6837\ : Span12Mux_s9_v
    port map (
            O => \N__34993\,
            I => \N__34987\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__34990\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6835\ : Odrv12
    port map (
            O => \N__34987\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6834\ : CascadeMux
    port map (
            O => \N__34982\,
            I => \N__34979\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34976\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__34976\,
            I => \N__34972\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34969\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__34972\,
            I => \N__34966\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34963\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__34966\,
            I => \N__34955\
        );

    \I__6827\ : Span4Mux_v
    port map (
            O => \N__34963\,
            I => \N__34955\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34948\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34948\
        );

    \I__6824\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34948\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__34955\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__34948\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34938\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34935\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__34941\,
            I => \N__34932\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__34938\,
            I => \N__34929\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34935\,
            I => \N__34926\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34922\
        );

    \I__6815\ : Span4Mux_v
    port map (
            O => \N__34929\,
            I => \N__34919\
        );

    \I__6814\ : Span12Mux_v
    port map (
            O => \N__34926\,
            I => \N__34916\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34913\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34922\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6811\ : Odrv4
    port map (
            O => \N__34919\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6810\ : Odrv12
    port map (
            O => \N__34916\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__34913\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6808\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34899\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34894\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34894\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__34899\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34894\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__34889\,
            I => \N__34885\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__34888\,
            I => \N__34881\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34878\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34875\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34872\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34878\,
            I => \N__34869\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34875\,
            I => \N__34864\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__34872\,
            I => \N__34864\
        );

    \I__6795\ : Span12Mux_h
    port map (
            O => \N__34869\,
            I => \N__34861\
        );

    \I__6794\ : Span12Mux_v
    port map (
            O => \N__34864\,
            I => \N__34858\
        );

    \I__6793\ : Span12Mux_v
    port map (
            O => \N__34861\,
            I => \N__34855\
        );

    \I__6792\ : Odrv12
    port map (
            O => \N__34858\,
            I => \il_min_comp1_D2\
        );

    \I__6791\ : Odrv12
    port map (
            O => \N__34855\,
            I => \il_min_comp1_D2\
        );

    \I__6790\ : CascadeMux
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34844\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__34844\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34838\,
            I => \N__34833\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34830\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34827\
        );

    \I__6783\ : Span4Mux_v
    port map (
            O => \N__34833\,
            I => \N__34824\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34830\,
            I => \N__34821\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34811\
        );

    \I__6780\ : Span4Mux_h
    port map (
            O => \N__34824\,
            I => \N__34811\
        );

    \I__6779\ : Span4Mux_h
    port map (
            O => \N__34821\,
            I => \N__34811\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34806\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34806\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34803\
        );

    \I__6775\ : Odrv4
    port map (
            O => \N__34811\,
            I => phase_controller_inst1_state_4
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__34806\,
            I => phase_controller_inst1_state_4
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__34803\,
            I => phase_controller_inst1_state_4
        );

    \I__6772\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34793\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__34793\,
            I => \N__34789\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34786\
        );

    \I__6769\ : Odrv4
    port map (
            O => \N__34789\,
            I => \phase_controller_inst1.N_54\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__34786\,
            I => \phase_controller_inst1.N_54\
        );

    \I__6767\ : CascadeMux
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34778\,
            I => \N__34775\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__34775\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34769\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__34769\,
            I => \N__34764\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34761\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34758\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__34764\,
            I => \N__34755\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__34761\,
            I => \N__34752\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__34758\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__6757\ : Odrv4
    port map (
            O => \N__34755\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__6756\ : Odrv12
    port map (
            O => \N__34752\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34740\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34744\,
            I => \N__34737\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34734\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34740\,
            I => \N__34731\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34737\,
            I => \N__34728\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__34734\,
            I => \N__34725\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__34731\,
            I => \N__34721\
        );

    \I__6748\ : Span4Mux_v
    port map (
            O => \N__34728\,
            I => \N__34716\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__34725\,
            I => \N__34716\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34713\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__34721\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__34716\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__34713\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__34706\,
            I => \N__34690\
        );

    \I__6741\ : CascadeMux
    port map (
            O => \N__34705\,
            I => \N__34669\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34651\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34651\
        );

    \I__6738\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34651\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34651\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34651\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34642\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34642\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34642\
        );

    \I__6732\ : InMux
    port map (
            O => \N__34696\,
            I => \N__34642\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34629\
        );

    \I__6730\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34629\
        );

    \I__6729\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34629\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34690\,
            I => \N__34629\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34689\,
            I => \N__34629\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34629\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34687\,
            I => \N__34626\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34617\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34617\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__34684\,
            I => \N__34599\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34579\
        );

    \I__6720\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34579\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34579\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34562\
        );

    \I__6717\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34562\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34562\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34562\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34562\
        );

    \I__6713\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34562\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34674\,
            I => \N__34551\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34551\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34551\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34669\,
            I => \N__34551\
        );

    \I__6708\ : InMux
    port map (
            O => \N__34668\,
            I => \N__34551\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34538\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34666\,
            I => \N__34538\
        );

    \I__6705\ : InMux
    port map (
            O => \N__34665\,
            I => \N__34538\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34538\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34663\,
            I => \N__34538\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34538\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__34651\,
            I => \N__34533\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__34642\,
            I => \N__34533\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__34629\,
            I => \N__34529\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__34626\,
            I => \N__34526\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34521\
        );

    \I__6696\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34521\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34516\
        );

    \I__6694\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34516\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__34617\,
            I => \N__34508\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34501\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34615\,
            I => \N__34501\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34501\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34496\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34496\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34491\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34491\
        );

    \I__6685\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34488\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34485\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__34607\,
            I => \N__34477\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34473\
        );

    \I__6681\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34457\
        );

    \I__6680\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34457\
        );

    \I__6679\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34457\
        );

    \I__6678\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34457\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34457\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34454\
        );

    \I__6675\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34441\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34596\,
            I => \N__34441\
        );

    \I__6673\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34441\
        );

    \I__6672\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34441\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34441\
        );

    \I__6670\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34441\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34430\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34430\
        );

    \I__6667\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34430\
        );

    \I__6666\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34430\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34430\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34586\,
            I => \N__34427\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__34579\,
            I => \N__34424\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34415\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34415\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34415\
        );

    \I__6659\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34415\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__34562\,
            I => \N__34406\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__34551\,
            I => \N__34406\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34406\
        );

    \I__6655\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34406\
        );

    \I__6654\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34403\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__34529\,
            I => \N__34396\
        );

    \I__6652\ : Span4Mux_v
    port map (
            O => \N__34526\,
            I => \N__34396\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__34521\,
            I => \N__34396\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__34516\,
            I => \N__34393\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34382\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34382\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34382\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34382\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34382\
        );

    \I__6644\ : Span4Mux_v
    port map (
            O => \N__34508\,
            I => \N__34377\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__34501\,
            I => \N__34377\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34372\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__34491\,
            I => \N__34372\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__34488\,
            I => \N__34369\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34485\,
            I => \N__34366\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34359\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34359\
        );

    \I__6636\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34359\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34354\
        );

    \I__6634\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34354\
        );

    \I__6633\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34349\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34349\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34346\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34335\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34335\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34335\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34335\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34335\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__34457\,
            I => \N__34326\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__34454\,
            I => \N__34326\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34326\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__34430\,
            I => \N__34326\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__34427\,
            I => \N__34317\
        );

    \I__6620\ : Span4Mux_v
    port map (
            O => \N__34424\,
            I => \N__34317\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__34415\,
            I => \N__34317\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__34406\,
            I => \N__34317\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34312\
        );

    \I__6616\ : Span4Mux_h
    port map (
            O => \N__34396\,
            I => \N__34312\
        );

    \I__6615\ : Span4Mux_h
    port map (
            O => \N__34393\,
            I => \N__34301\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34301\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__34377\,
            I => \N__34301\
        );

    \I__6612\ : Span4Mux_h
    port map (
            O => \N__34372\,
            I => \N__34301\
        );

    \I__6611\ : Span4Mux_h
    port map (
            O => \N__34369\,
            I => \N__34301\
        );

    \I__6610\ : Span12Mux_s10_h
    port map (
            O => \N__34366\,
            I => \N__34298\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__34359\,
            I => \N__34291\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__34354\,
            I => \N__34291\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34291\
        );

    \I__6606\ : Odrv4
    port map (
            O => \N__34346\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__34335\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6604\ : Odrv12
    port map (
            O => \N__34326\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__34317\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__34312\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6601\ : Odrv4
    port map (
            O => \N__34301\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6600\ : Odrv12
    port map (
            O => \N__34298\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__34291\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__34274\,
            I => \N__34270\
        );

    \I__6597\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34265\
        );

    \I__6596\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34265\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__34265\,
            I => \N__34262\
        );

    \I__6594\ : Odrv12
    port map (
            O => \N__34262\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__6593\ : CEMux
    port map (
            O => \N__34259\,
            I => \N__34255\
        );

    \I__6592\ : CEMux
    port map (
            O => \N__34258\,
            I => \N__34239\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34236\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34229\
        );

    \I__6589\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34229\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34252\,
            I => \N__34229\
        );

    \I__6587\ : CEMux
    port map (
            O => \N__34251\,
            I => \N__34226\
        );

    \I__6586\ : CEMux
    port map (
            O => \N__34250\,
            I => \N__34223\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34214\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34214\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34214\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34214\
        );

    \I__6581\ : CEMux
    port map (
            O => \N__34245\,
            I => \N__34211\
        );

    \I__6580\ : CEMux
    port map (
            O => \N__34244\,
            I => \N__34208\
        );

    \I__6579\ : CEMux
    port map (
            O => \N__34243\,
            I => \N__34196\
        );

    \I__6578\ : CEMux
    port map (
            O => \N__34242\,
            I => \N__34193\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__34239\,
            I => \N__34186\
        );

    \I__6576\ : Span4Mux_h
    port map (
            O => \N__34236\,
            I => \N__34170\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34229\,
            I => \N__34170\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__34226\,
            I => \N__34167\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34156\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__34214\,
            I => \N__34156\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34211\,
            I => \N__34156\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34152\
        );

    \I__6569\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34145\
        );

    \I__6568\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34145\
        );

    \I__6567\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34145\
        );

    \I__6566\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34134\
        );

    \I__6565\ : InMux
    port map (
            O => \N__34203\,
            I => \N__34134\
        );

    \I__6564\ : InMux
    port map (
            O => \N__34202\,
            I => \N__34134\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34134\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34134\
        );

    \I__6561\ : CEMux
    port map (
            O => \N__34199\,
            I => \N__34131\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__34196\,
            I => \N__34128\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__34193\,
            I => \N__34125\
        );

    \I__6558\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34116\
        );

    \I__6557\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34116\
        );

    \I__6556\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34116\
        );

    \I__6555\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34116\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__34186\,
            I => \N__34113\
        );

    \I__6553\ : CEMux
    port map (
            O => \N__34185\,
            I => \N__34110\
        );

    \I__6552\ : CEMux
    port map (
            O => \N__34184\,
            I => \N__34107\
        );

    \I__6551\ : CEMux
    port map (
            O => \N__34183\,
            I => \N__34104\
        );

    \I__6550\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34095\
        );

    \I__6549\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34095\
        );

    \I__6548\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34095\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34095\
        );

    \I__6546\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34086\
        );

    \I__6545\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34086\
        );

    \I__6544\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34086\
        );

    \I__6543\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34086\
        );

    \I__6542\ : Span4Mux_v
    port map (
            O => \N__34170\,
            I => \N__34081\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__34167\,
            I => \N__34081\
        );

    \I__6540\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34072\
        );

    \I__6539\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34072\
        );

    \I__6538\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34072\
        );

    \I__6537\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34072\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__34156\,
            I => \N__34069\
        );

    \I__6535\ : CEMux
    port map (
            O => \N__34155\,
            I => \N__34066\
        );

    \I__6534\ : Span4Mux_h
    port map (
            O => \N__34152\,
            I => \N__34063\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34145\,
            I => \N__34058\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__34134\,
            I => \N__34058\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__34131\,
            I => \N__34055\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__34128\,
            I => \N__34052\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__34125\,
            I => \N__34049\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__34116\,
            I => \N__34046\
        );

    \I__6527\ : Span4Mux_v
    port map (
            O => \N__34113\,
            I => \N__34039\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__34110\,
            I => \N__34039\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__34107\,
            I => \N__34039\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__34104\,
            I => \N__34032\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__34095\,
            I => \N__34032\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__34086\,
            I => \N__34032\
        );

    \I__6521\ : Span4Mux_h
    port map (
            O => \N__34081\,
            I => \N__34025\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__34072\,
            I => \N__34025\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__34069\,
            I => \N__34025\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__34066\,
            I => \N__34018\
        );

    \I__6517\ : Span4Mux_h
    port map (
            O => \N__34063\,
            I => \N__34018\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__34058\,
            I => \N__34018\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__34055\,
            I => \N__34009\
        );

    \I__6514\ : Span4Mux_h
    port map (
            O => \N__34052\,
            I => \N__34009\
        );

    \I__6513\ : Span4Mux_h
    port map (
            O => \N__34049\,
            I => \N__34009\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__34046\,
            I => \N__34009\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__34039\,
            I => \N__34006\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__34032\,
            I => \N__34001\
        );

    \I__6509\ : Span4Mux_v
    port map (
            O => \N__34025\,
            I => \N__34001\
        );

    \I__6508\ : Span4Mux_v
    port map (
            O => \N__34018\,
            I => \N__33998\
        );

    \I__6507\ : Span4Mux_v
    port map (
            O => \N__34009\,
            I => \N__33995\
        );

    \I__6506\ : Odrv4
    port map (
            O => \N__34006\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__34001\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__33998\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__33995\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33983\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__33983\,
            I => \N__33979\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33976\
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__33979\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__33976\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33968\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33968\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33961\
        );

    \I__6494\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33958\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33955\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33958\,
            I => \N__33952\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__33955\,
            I => \N__33948\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__33952\,
            I => \N__33945\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33942\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__33948\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33945\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33942\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6485\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33932\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__33932\,
            I => \N__33929\
        );

    \I__6483\ : Span4Mux_v
    port map (
            O => \N__33929\,
            I => \N__33926\
        );

    \I__6482\ : Odrv4
    port map (
            O => \N__33926\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__6481\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33919\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33916\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33919\,
            I => \N__33913\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33916\,
            I => \N__33909\
        );

    \I__6477\ : Span4Mux_h
    port map (
            O => \N__33913\,
            I => \N__33906\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33903\
        );

    \I__6475\ : Odrv12
    port map (
            O => \N__33909\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__6474\ : Odrv4
    port map (
            O => \N__33906\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__33903\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__6472\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33893\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33893\,
            I => \N__33890\
        );

    \I__6470\ : Odrv12
    port map (
            O => \N__33890\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33883\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__33886\,
            I => \N__33880\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33874\
        );

    \I__6465\ : Span4Mux_h
    port map (
            O => \N__33877\,
            I => \N__33871\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33868\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__33871\,
            I => \N__33864\
        );

    \I__6462\ : Span4Mux_h
    port map (
            O => \N__33868\,
            I => \N__33861\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33867\,
            I => \N__33858\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__33864\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6459\ : Odrv4
    port map (
            O => \N__33861\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__33858\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33845\
        );

    \I__6455\ : Odrv12
    port map (
            O => \N__33845\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33839\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__33839\,
            I => \N__33835\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33832\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__33835\,
            I => \N__33829\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__33832\,
            I => \N__33826\
        );

    \I__6449\ : Span4Mux_h
    port map (
            O => \N__33829\,
            I => \N__33820\
        );

    \I__6448\ : Span4Mux_v
    port map (
            O => \N__33826\,
            I => \N__33820\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33817\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__33820\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__33817\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33809\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33809\,
            I => \N__33806\
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__33806\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33800\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33794\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33794\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__6437\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33788\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__33782\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33776\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__33776\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33770\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33770\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33764\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__33764\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33758\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__33758\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33752\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33752\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__6423\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33746\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33743\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__33743\,
            I => \N__33740\
        );

    \I__6420\ : Sp12to4
    port map (
            O => \N__33740\,
            I => \N__33737\
        );

    \I__6419\ : Span12Mux_v
    port map (
            O => \N__33737\,
            I => \N__33734\
        );

    \I__6418\ : Odrv12
    port map (
            O => \N__33734\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33728\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__33728\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__6415\ : CascadeMux
    port map (
            O => \N__33725\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33719\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__33716\,
            I => \N__33712\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33709\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__33712\,
            I => \N__33706\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33703\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__33706\,
            I => \N__33700\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__33703\,
            I => \N__33697\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__33700\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__33697\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__33692\,
            I => \N__33687\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33684\
        );

    \I__6402\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33681\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33678\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__33684\,
            I => \current_shift_inst.N_1326_i\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33681\,
            I => \current_shift_inst.N_1326_i\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__33678\,
            I => \current_shift_inst.N_1326_i\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33665\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__33665\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__6394\ : CascadeMux
    port map (
            O => \N__33662\,
            I => \phase_controller_inst1.N_55_cascade_\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33656\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33656\,
            I => \N__33653\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__33653\,
            I => \N__33649\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33646\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__33649\,
            I => state_ns_i_a2_1
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33646\,
            I => state_ns_i_a2_1
        );

    \I__6387\ : InMux
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33633\
        );

    \I__6385\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33630\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33627\
        );

    \I__6383\ : Span4Mux_v
    port map (
            O => \N__33633\,
            I => \N__33622\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33622\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__33627\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__33622\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6379\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__33614\,
            I => \N__33611\
        );

    \I__6377\ : Span4Mux_v
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__6376\ : Span4Mux_h
    port map (
            O => \N__33608\,
            I => \N__33605\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__33605\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__6374\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33599\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__33599\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__6372\ : IoInMux
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33593\,
            I => \N__33590\
        );

    \I__6370\ : Span4Mux_s2_v
    port map (
            O => \N__33590\,
            I => \N__33587\
        );

    \I__6369\ : Sp12to4
    port map (
            O => \N__33587\,
            I => \N__33584\
        );

    \I__6368\ : Span12Mux_h
    port map (
            O => \N__33584\,
            I => \N__33580\
        );

    \I__6367\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33577\
        );

    \I__6366\ : Odrv12
    port map (
            O => \N__33580\,
            I => \T23_c\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33577\,
            I => \T23_c\
        );

    \I__6364\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33566\
        );

    \I__6363\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33566\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__33566\,
            I => \N__33561\
        );

    \I__6361\ : InMux
    port map (
            O => \N__33565\,
            I => \N__33556\
        );

    \I__6360\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33556\
        );

    \I__6359\ : Odrv12
    port map (
            O => \N__33561\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__33556\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6357\ : IoInMux
    port map (
            O => \N__33551\,
            I => \N__33548\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33545\
        );

    \I__6355\ : IoSpan4Mux
    port map (
            O => \N__33545\,
            I => \N__33542\
        );

    \I__6354\ : Span4Mux_s3_v
    port map (
            O => \N__33542\,
            I => \N__33539\
        );

    \I__6353\ : Span4Mux_v
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__6352\ : Span4Mux_v
    port map (
            O => \N__33536\,
            I => \N__33532\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33529\
        );

    \I__6350\ : Odrv4
    port map (
            O => \N__33532\,
            I => \T45_c\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__33529\,
            I => \T45_c\
        );

    \I__6348\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33520\
        );

    \I__6347\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33517\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__33520\,
            I => \N__33514\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__33517\,
            I => \N__33511\
        );

    \I__6344\ : Span4Mux_h
    port map (
            O => \N__33514\,
            I => \N__33508\
        );

    \I__6343\ : Span12Mux_v
    port map (
            O => \N__33511\,
            I => \N__33504\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__33508\,
            I => \N__33501\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33498\
        );

    \I__6340\ : Odrv12
    port map (
            O => \N__33504\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__6339\ : Odrv4
    port map (
            O => \N__33501\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33498\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__6335\ : Odrv4
    port map (
            O => \N__33485\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__33482\,
            I => \N__33478\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33481\,
            I => \N__33475\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33472\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33475\,
            I => \N__33469\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__33472\,
            I => \N__33466\
        );

    \I__6329\ : Span4Mux_v
    port map (
            O => \N__33469\,
            I => \N__33462\
        );

    \I__6328\ : Span4Mux_h
    port map (
            O => \N__33466\,
            I => \N__33459\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33456\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__33462\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6325\ : Odrv4
    port map (
            O => \N__33459\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__33456\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33443\
        );

    \I__6321\ : Odrv4
    port map (
            O => \N__33443\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__6320\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33436\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33433\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33427\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__33433\,
            I => \N__33427\
        );

    \I__6316\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33424\
        );

    \I__6315\ : Span4Mux_h
    port map (
            O => \N__33427\,
            I => \N__33421\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__33424\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__6313\ : Odrv4
    port map (
            O => \N__33421\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__33416\,
            I => \N__33413\
        );

    \I__6311\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33409\
        );

    \I__6310\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33406\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__33409\,
            I => \N__33400\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__33406\,
            I => \N__33400\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33397\
        );

    \I__6306\ : Span4Mux_h
    port map (
            O => \N__33400\,
            I => \N__33394\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__33397\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__6304\ : Odrv4
    port map (
            O => \N__33394\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__6303\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33385\
        );

    \I__6302\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33382\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33379\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__33382\,
            I => \N__33376\
        );

    \I__6299\ : Span4Mux_v
    port map (
            O => \N__33379\,
            I => \N__33373\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__33376\,
            I => \N__33369\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__33373\,
            I => \N__33366\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33363\
        );

    \I__6295\ : Odrv4
    port map (
            O => \N__33369\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6294\ : Odrv4
    port map (
            O => \N__33366\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__33363\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33353\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33350\
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__33350\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__6289\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33344\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__33344\,
            I => \N__33339\
        );

    \I__6287\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33336\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33342\,
            I => \N__33333\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__33339\,
            I => \N__33328\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33336\,
            I => \N__33328\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__33333\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__33328\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33323\,
            I => \N__33320\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__33320\,
            I => \N__33315\
        );

    \I__6279\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33312\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33309\
        );

    \I__6277\ : Span4Mux_v
    port map (
            O => \N__33315\,
            I => \N__33304\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__33312\,
            I => \N__33304\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__33309\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6274\ : Odrv4
    port map (
            O => \N__33304\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__33299\,
            I => \N__33295\
        );

    \I__6272\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33292\
        );

    \I__6271\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33289\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__33292\,
            I => \N__33286\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__33289\,
            I => \N__33283\
        );

    \I__6268\ : Span4Mux_h
    port map (
            O => \N__33286\,
            I => \N__33279\
        );

    \I__6267\ : Span4Mux_v
    port map (
            O => \N__33283\,
            I => \N__33276\
        );

    \I__6266\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33273\
        );

    \I__6265\ : Odrv4
    port map (
            O => \N__33279\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__33276\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__33273\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6262\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33263\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__33263\,
            I => \N__33260\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__33260\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33254\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33251\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__33251\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33248\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33242\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33239\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__33239\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33236\,
            I => \bfn_12_14_0_\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33230\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__33230\,
            I => \N__33227\
        );

    \I__6249\ : Odrv12
    port map (
            O => \N__33227\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__6248\ : InMux
    port map (
            O => \N__33224\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33218\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__33218\,
            I => \N__33215\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__33215\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__6244\ : InMux
    port map (
            O => \N__33212\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__6243\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__33203\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__6240\ : InMux
    port map (
            O => \N__33200\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__6239\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33194\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33191\
        );

    \I__6237\ : Odrv12
    port map (
            O => \N__33191\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__6236\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33181\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33181\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33178\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33181\,
            I => \N__33175\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__33178\,
            I => \N__33172\
        );

    \I__6231\ : Span4Mux_h
    port map (
            O => \N__33175\,
            I => \N__33169\
        );

    \I__6230\ : Odrv12
    port map (
            O => \N__33172\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__33169\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33164\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__6227\ : InMux
    port map (
            O => \N__33161\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33158\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__33152\,
            I => \N__33148\
        );

    \I__6223\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33145\
        );

    \I__6222\ : Span4Mux_h
    port map (
            O => \N__33148\,
            I => \N__33142\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__33145\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__33142\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33134\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__33134\,
            I => \N__33131\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__33131\,
            I => \N__33128\
        );

    \I__6216\ : Span4Mux_h
    port map (
            O => \N__33128\,
            I => \N__33125\
        );

    \I__6215\ : Odrv4
    port map (
            O => \N__33125\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33119\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__33119\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__6212\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33113\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__33113\,
            I => \N__33110\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__33110\,
            I => \current_shift_inst.control_input_18\
        );

    \I__6209\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33104\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__33104\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__6207\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33098\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__33098\,
            I => \N__33095\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__33095\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__6204\ : InMux
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__33089\,
            I => \N__33085\
        );

    \I__6202\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33082\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__33085\,
            I => \N__33077\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__33082\,
            I => \N__33077\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__33077\,
            I => \N__33074\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__33074\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6197\ : InMux
    port map (
            O => \N__33071\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__33068\,
            I => \N__33065\
        );

    \I__6195\ : InMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33059\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__33059\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__6192\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33053\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__33053\,
            I => \N__33049\
        );

    \I__6190\ : InMux
    port map (
            O => \N__33052\,
            I => \N__33046\
        );

    \I__6189\ : Span4Mux_h
    port map (
            O => \N__33049\,
            I => \N__33041\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__33046\,
            I => \N__33041\
        );

    \I__6187\ : Span4Mux_h
    port map (
            O => \N__33041\,
            I => \N__33038\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__33038\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6185\ : InMux
    port map (
            O => \N__33035\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__6184\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__33029\,
            I => \N__33026\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__33026\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__6181\ : InMux
    port map (
            O => \N__33023\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__6180\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33017\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__33017\,
            I => \N__33014\
        );

    \I__6178\ : Odrv12
    port map (
            O => \N__33014\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__6177\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33008\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__33008\,
            I => \N__33003\
        );

    \I__6175\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32998\
        );

    \I__6174\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32998\
        );

    \I__6173\ : Span4Mux_v
    port map (
            O => \N__33003\,
            I => \N__32995\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__32998\,
            I => \N__32992\
        );

    \I__6171\ : Span4Mux_h
    port map (
            O => \N__32995\,
            I => \N__32987\
        );

    \I__6170\ : Span4Mux_v
    port map (
            O => \N__32992\,
            I => \N__32987\
        );

    \I__6169\ : Odrv4
    port map (
            O => \N__32987\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32984\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32978\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32975\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__32975\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32972\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32966\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__32966\,
            I => \N__32963\
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__32963\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__6160\ : InMux
    port map (
            O => \N__32960\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32957\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__6158\ : InMux
    port map (
            O => \N__32954\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32951\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32948\,
            I => \bfn_12_12_0_\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32945\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32942\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32939\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__6152\ : InMux
    port map (
            O => \N__32936\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32933\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__32930\,
            I => \N__32926\
        );

    \I__6149\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32923\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32918\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__32923\,
            I => \N__32915\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__32922\,
            I => \N__32912\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32909\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32918\,
            I => \N__32906\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__32915\,
            I => \N__32903\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32900\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32909\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6140\ : Odrv12
    port map (
            O => \N__32906\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6139\ : Odrv4
    port map (
            O => \N__32903\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32900\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32884\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32887\,
            I => \N__32880\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__32884\,
            I => \N__32877\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32874\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32880\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__32877\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__32874\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32863\
        );

    \I__6128\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32860\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32863\,
            I => \N__32857\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__32860\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__6125\ : Odrv12
    port map (
            O => \N__32857\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__32852\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32843\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32843\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32839\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32835\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__32839\,
            I => \N__32832\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32829\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32835\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__32832\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__32829\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6114\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32819\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32816\
        );

    \I__6112\ : Span4Mux_v
    port map (
            O => \N__32816\,
            I => \N__32813\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__32813\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32806\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32801\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32806\,
            I => \N__32798\
        );

    \I__6107\ : CascadeMux
    port map (
            O => \N__32805\,
            I => \N__32795\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32792\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32787\
        );

    \I__6104\ : Span4Mux_v
    port map (
            O => \N__32798\,
            I => \N__32787\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32784\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__32792\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6101\ : Odrv4
    port map (
            O => \N__32787\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32784\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6099\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32774\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__32774\,
            I => \N__32770\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32773\,
            I => \N__32766\
        );

    \I__6096\ : Span4Mux_h
    port map (
            O => \N__32770\,
            I => \N__32763\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32760\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__32766\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__32763\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__32760\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32753\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__6090\ : InMux
    port map (
            O => \N__32750\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32747\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32744\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32738\,
            I => \il_min_comp1_D1\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32732\,
            I => \N__32727\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32724\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32721\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__32727\,
            I => \N__32718\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32713\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__32721\,
            I => \N__32713\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__32718\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__6077\ : Odrv12
    port map (
            O => \N__32713\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32704\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32701\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32704\,
            I => \N__32696\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__32701\,
            I => \N__32693\
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__32700\,
            I => \N__32690\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32699\,
            I => \N__32687\
        );

    \I__6070\ : Span4Mux_h
    port map (
            O => \N__32696\,
            I => \N__32682\
        );

    \I__6069\ : Span4Mux_h
    port map (
            O => \N__32693\,
            I => \N__32682\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32679\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32687\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__32682\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32679\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32666\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32666\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__32666\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32659\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32655\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32659\,
            I => \N__32652\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32649\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__32655\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__6056\ : Odrv12
    port map (
            O => \N__32652\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32649\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__6054\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32639\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32639\,
            I => \N__32635\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32631\
        );

    \I__6051\ : Span4Mux_h
    port map (
            O => \N__32635\,
            I => \N__32627\
        );

    \I__6050\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32624\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__32631\,
            I => \N__32621\
        );

    \I__6048\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32618\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__32627\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__32624\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__6045\ : Odrv12
    port map (
            O => \N__32621\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__32618\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__6043\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32606\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32603\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__32603\,
            I => \N__32600\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__32600\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32594\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__32594\,
            I => \N__32591\
        );

    \I__6037\ : Span4Mux_v
    port map (
            O => \N__32591\,
            I => \N__32588\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__32588\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__6035\ : CascadeMux
    port map (
            O => \N__32585\,
            I => \N__32581\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32584\,
            I => \N__32577\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32574\
        );

    \I__6032\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32571\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__32577\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__32574\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32571\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6028\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32559\
        );

    \I__6027\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32554\
        );

    \I__6026\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32554\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32559\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32554\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__32549\,
            I => \N__32545\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32540\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32540\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__32540\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__6019\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32533\
        );

    \I__6018\ : InMux
    port map (
            O => \N__32536\,
            I => \N__32530\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__32533\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__32530\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__32525\,
            I => \N__32522\
        );

    \I__6014\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32519\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__32519\,
            I => \N__32516\
        );

    \I__6012\ : Span4Mux_v
    port map (
            O => \N__32516\,
            I => \N__32513\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__32513\,
            I => \N__32510\
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__32510\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32500\
        );

    \I__6007\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32496\
        );

    \I__6006\ : Span4Mux_h
    port map (
            O => \N__32500\,
            I => \N__32493\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32490\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__32496\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__32493\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__32490\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32480\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__32480\,
            I => \N__32476\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32472\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__32476\,
            I => \N__32469\
        );

    \I__5997\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32466\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__32472\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__32469\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__5993\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32456\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__32456\,
            I => \N__32452\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32448\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__32452\,
            I => \N__32445\
        );

    \I__5989\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32442\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__32448\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__32445\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__32442\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__32435\,
            I => \N__32432\
        );

    \I__5984\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32429\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32429\,
            I => \N__32425\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32421\
        );

    \I__5981\ : Span4Mux_h
    port map (
            O => \N__32425\,
            I => \N__32418\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32415\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__32421\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5978\ : Odrv4
    port map (
            O => \N__32418\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__32415\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32405\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32402\
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__32402\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__32399\,
            I => \N__32376\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__32398\,
            I => \N__32373\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32370\
        );

    \I__5970\ : CascadeMux
    port map (
            O => \N__32396\,
            I => \N__32362\
        );

    \I__5969\ : CascadeMux
    port map (
            O => \N__32395\,
            I => \N__32359\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__32394\,
            I => \N__32356\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__32393\,
            I => \N__32353\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32343\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32343\
        );

    \I__5964\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32343\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32332\
        );

    \I__5962\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32332\
        );

    \I__5961\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32332\
        );

    \I__5960\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32332\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32332\
        );

    \I__5958\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32329\
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__32383\,
            I => \N__32323\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__32382\,
            I => \N__32320\
        );

    \I__5955\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32309\
        );

    \I__5954\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32309\
        );

    \I__5953\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32309\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32309\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32309\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__32370\,
            I => \N__32306\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32299\
        );

    \I__5948\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32299\
        );

    \I__5947\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32299\
        );

    \I__5946\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32292\
        );

    \I__5945\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32292\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32292\
        );

    \I__5943\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32279\
        );

    \I__5942\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32279\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32279\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32279\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32279\
        );

    \I__5938\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32279\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32276\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__32332\,
            I => \N__32273\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__32329\,
            I => \N__32270\
        );

    \I__5934\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32259\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32259\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32259\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32259\
        );

    \I__5930\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32259\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32254\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__32306\,
            I => \N__32254\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32249\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32292\,
            I => \N__32249\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32246\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__32276\,
            I => \N__32241\
        );

    \I__5923\ : Span4Mux_v
    port map (
            O => \N__32273\,
            I => \N__32241\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__32270\,
            I => \N__32238\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32259\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__32254\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__5919\ : Odrv12
    port map (
            O => \N__32249\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__32246\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__32241\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__32238\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__32225\,
            I => \N__32220\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__32224\,
            I => \N__32216\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__32223\,
            I => \N__32208\
        );

    \I__5912\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32205\
        );

    \I__5911\ : CascadeMux
    port map (
            O => \N__32219\,
            I => \N__32194\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32189\
        );

    \I__5909\ : CascadeMux
    port map (
            O => \N__32215\,
            I => \N__32184\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__32214\,
            I => \N__32181\
        );

    \I__5907\ : CascadeMux
    port map (
            O => \N__32213\,
            I => \N__32178\
        );

    \I__5906\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32171\
        );

    \I__5905\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32171\
        );

    \I__5904\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32171\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32168\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__32204\,
            I => \N__32165\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__32203\,
            I => \N__32162\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__32202\,
            I => \N__32159\
        );

    \I__5899\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32142\
        );

    \I__5898\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32142\
        );

    \I__5897\ : InMux
    port map (
            O => \N__32199\,
            I => \N__32142\
        );

    \I__5896\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32142\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32142\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32135\
        );

    \I__5893\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32135\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32192\,
            I => \N__32135\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__32189\,
            I => \N__32127\
        );

    \I__5890\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32116\
        );

    \I__5889\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32116\
        );

    \I__5888\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32116\
        );

    \I__5887\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32116\
        );

    \I__5886\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32116\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__32171\,
            I => \N__32113\
        );

    \I__5884\ : Span4Mux_v
    port map (
            O => \N__32168\,
            I => \N__32110\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32103\
        );

    \I__5882\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32103\
        );

    \I__5881\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32103\
        );

    \I__5880\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32096\
        );

    \I__5879\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32096\
        );

    \I__5878\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32096\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32089\
        );

    \I__5876\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32089\
        );

    \I__5875\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32089\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__32142\,
            I => \N__32084\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__32135\,
            I => \N__32084\
        );

    \I__5872\ : InMux
    port map (
            O => \N__32134\,
            I => \N__32073\
        );

    \I__5871\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32073\
        );

    \I__5870\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32073\
        );

    \I__5869\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32073\
        );

    \I__5868\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32073\
        );

    \I__5867\ : Sp12to4
    port map (
            O => \N__32127\,
            I => \N__32068\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__32116\,
            I => \N__32068\
        );

    \I__5865\ : Span4Mux_h
    port map (
            O => \N__32113\,
            I => \N__32065\
        );

    \I__5864\ : Sp12to4
    port map (
            O => \N__32110\,
            I => \N__32056\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32056\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32056\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32056\
        );

    \I__5860\ : Span4Mux_v
    port map (
            O => \N__32084\,
            I => \N__32053\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32048\
        );

    \I__5858\ : Span12Mux_v
    port map (
            O => \N__32068\,
            I => \N__32048\
        );

    \I__5857\ : Span4Mux_v
    port map (
            O => \N__32065\,
            I => \N__32045\
        );

    \I__5856\ : Span12Mux_h
    port map (
            O => \N__32056\,
            I => \N__32042\
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__32053\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__5854\ : Odrv12
    port map (
            O => \N__32048\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__5853\ : Odrv4
    port map (
            O => \N__32045\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__5852\ : Odrv12
    port map (
            O => \N__32042\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__5851\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32010\
        );

    \I__5850\ : InMux
    port map (
            O => \N__32032\,
            I => \N__32006\
        );

    \I__5849\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32000\
        );

    \I__5848\ : InMux
    port map (
            O => \N__32030\,
            I => \N__31993\
        );

    \I__5847\ : InMux
    port map (
            O => \N__32029\,
            I => \N__31993\
        );

    \I__5846\ : InMux
    port map (
            O => \N__32028\,
            I => \N__31993\
        );

    \I__5845\ : InMux
    port map (
            O => \N__32027\,
            I => \N__31981\
        );

    \I__5844\ : InMux
    port map (
            O => \N__32026\,
            I => \N__31981\
        );

    \I__5843\ : InMux
    port map (
            O => \N__32025\,
            I => \N__31981\
        );

    \I__5842\ : InMux
    port map (
            O => \N__32024\,
            I => \N__31981\
        );

    \I__5841\ : InMux
    port map (
            O => \N__32023\,
            I => \N__31981\
        );

    \I__5840\ : InMux
    port map (
            O => \N__32022\,
            I => \N__31970\
        );

    \I__5839\ : InMux
    port map (
            O => \N__32021\,
            I => \N__31970\
        );

    \I__5838\ : InMux
    port map (
            O => \N__32020\,
            I => \N__31970\
        );

    \I__5837\ : InMux
    port map (
            O => \N__32019\,
            I => \N__31970\
        );

    \I__5836\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31970\
        );

    \I__5835\ : InMux
    port map (
            O => \N__32017\,
            I => \N__31959\
        );

    \I__5834\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31959\
        );

    \I__5833\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31959\
        );

    \I__5832\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31959\
        );

    \I__5831\ : InMux
    port map (
            O => \N__32013\,
            I => \N__31959\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__32010\,
            I => \N__31956\
        );

    \I__5829\ : InMux
    port map (
            O => \N__32009\,
            I => \N__31953\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__32006\,
            I => \N__31950\
        );

    \I__5827\ : InMux
    port map (
            O => \N__32005\,
            I => \N__31938\
        );

    \I__5826\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31938\
        );

    \I__5825\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31938\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__32000\,
            I => \N__31935\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31993\,
            I => \N__31932\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31929\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__31981\,
            I => \N__31926\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__31970\,
            I => \N__31923\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__31959\,
            I => \N__31919\
        );

    \I__5818\ : Span4Mux_v
    port map (
            O => \N__31956\,
            I => \N__31912\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31953\,
            I => \N__31912\
        );

    \I__5816\ : Span4Mux_v
    port map (
            O => \N__31950\,
            I => \N__31912\
        );

    \I__5815\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31901\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31901\
        );

    \I__5813\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31901\
        );

    \I__5812\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31901\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31901\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__31938\,
            I => \N__31894\
        );

    \I__5809\ : Span4Mux_v
    port map (
            O => \N__31935\,
            I => \N__31894\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__31932\,
            I => \N__31894\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31887\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__31926\,
            I => \N__31887\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__31923\,
            I => \N__31887\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31884\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__31919\,
            I => \N__31879\
        );

    \I__5802\ : Span4Mux_h
    port map (
            O => \N__31912\,
            I => \N__31879\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31901\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__31894\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__31887\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31884\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__31879\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__5796\ : CascadeMux
    port map (
            O => \N__31868\,
            I => \N__31865\
        );

    \I__5795\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31861\
        );

    \I__5794\ : CascadeMux
    port map (
            O => \N__31864\,
            I => \N__31858\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31861\,
            I => \N__31853\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31850\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31857\,
            I => \N__31847\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31856\,
            I => \N__31844\
        );

    \I__5789\ : Span4Mux_h
    port map (
            O => \N__31853\,
            I => \N__31838\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31850\,
            I => \N__31838\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__31847\,
            I => \N__31833\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31844\,
            I => \N__31833\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31830\
        );

    \I__5784\ : Span4Mux_h
    port map (
            O => \N__31838\,
            I => \N__31827\
        );

    \I__5783\ : Span12Mux_s11_h
    port map (
            O => \N__31833\,
            I => \N__31824\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31821\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__31827\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5780\ : Odrv12
    port map (
            O => \N__31824\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__31821\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__31808\,
            I => \N__31805\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__31805\,
            I => \N__31802\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__31802\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__31799\,
            I => \N__31791\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__31798\,
            I => \N__31787\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__31797\,
            I => \N__31783\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__31796\,
            I => \N__31779\
        );

    \I__5769\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31761\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31761\
        );

    \I__5767\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31761\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31761\
        );

    \I__5765\ : InMux
    port map (
            O => \N__31787\,
            I => \N__31761\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31761\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31761\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31761\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31752\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31752\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__31761\,
            I => \N__31749\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__31760\,
            I => \N__31746\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__31759\,
            I => \N__31742\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__31758\,
            I => \N__31738\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__31757\,
            I => \N__31734\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__31752\,
            I => \N__31730\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__31749\,
            I => \N__31727\
        );

    \I__5752\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31710\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31710\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31710\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31710\
        );

    \I__5748\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31710\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31710\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31710\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31710\
        );

    \I__5744\ : Span4Mux_h
    port map (
            O => \N__31730\,
            I => \N__31707\
        );

    \I__5743\ : Span4Mux_h
    port map (
            O => \N__31727\,
            I => \N__31704\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__31710\,
            I => \N__31701\
        );

    \I__5741\ : Span4Mux_h
    port map (
            O => \N__31707\,
            I => \N__31698\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__31704\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__5739\ : Odrv12
    port map (
            O => \N__31701\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__31698\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31688\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__31688\,
            I => \N__31685\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__31685\,
            I => \N__31682\
        );

    \I__5734\ : Span4Mux_v
    port map (
            O => \N__31682\,
            I => \N__31677\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31672\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31672\
        );

    \I__5731\ : Sp12to4
    port map (
            O => \N__31677\,
            I => \N__31667\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31672\,
            I => \N__31667\
        );

    \I__5729\ : Span12Mux_h
    port map (
            O => \N__31667\,
            I => \N__31664\
        );

    \I__5728\ : Span12Mux_v
    port map (
            O => \N__31664\,
            I => \N__31661\
        );

    \I__5727\ : Odrv12
    port map (
            O => \N__31661\,
            I => il_max_comp2_c
        );

    \I__5726\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31655\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31651\
        );

    \I__5724\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31646\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__31651\,
            I => \N__31643\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31650\,
            I => \N__31640\
        );

    \I__5721\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31637\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__31646\,
            I => \N__31634\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__31643\,
            I => \N__31631\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__31640\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__31637\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5716\ : Odrv12
    port map (
            O => \N__31634\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__31631\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5714\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__31619\,
            I => \N__31616\
        );

    \I__5712\ : Odrv4
    port map (
            O => \N__31616\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__31613\,
            I => \N__31610\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31607\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__31604\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__5707\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31598\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__31598\,
            I => \N__31595\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__31595\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__31592\,
            I => \N__31589\
        );

    \I__5703\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31586\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31583\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__31583\,
            I => \N__31580\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__31577\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31571\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31568\
        );

    \I__5696\ : Span4Mux_h
    port map (
            O => \N__31568\,
            I => \N__31565\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__31565\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__31562\,
            I => \N__31559\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31556\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__5690\ : Odrv4
    port map (
            O => \N__31550\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__5689\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__31541\,
            I => \N__31538\
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__31538\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__31535\,
            I => \N__31532\
        );

    \I__5684\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31528\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__31531\,
            I => \N__31525\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__31528\,
            I => \N__31522\
        );

    \I__5681\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31519\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__31522\,
            I => \N__31514\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__31519\,
            I => \N__31514\
        );

    \I__5678\ : Odrv4
    port map (
            O => \N__31514\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31508\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__31508\,
            I => \N__31505\
        );

    \I__5675\ : Sp12to4
    port map (
            O => \N__31505\,
            I => \N__31502\
        );

    \I__5674\ : Odrv12
    port map (
            O => \N__31502\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31499\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28\
        );

    \I__5672\ : InMux
    port map (
            O => \N__31496\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__5671\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31490\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__31490\,
            I => \N__31486\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31482\
        );

    \I__5668\ : Span4Mux_h
    port map (
            O => \N__31486\,
            I => \N__31479\
        );

    \I__5667\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31476\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31482\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__31479\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__31476\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__31469\,
            I => \N__31466\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31462\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31458\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__31462\,
            I => \N__31455\
        );

    \I__5659\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31452\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__31458\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__31455\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__31452\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5655\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31442\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__31442\,
            I => \N__31437\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \N__31434\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31440\,
            I => \N__31431\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__31437\,
            I => \N__31428\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31425\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__31431\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__31428\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__31425\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31415\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__31415\,
            I => \N__31411\
        );

    \I__5644\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31407\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__31411\,
            I => \N__31404\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31401\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__31407\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__31404\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__31401\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31388\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31385\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__31385\,
            I => \N__31382\
        );

    \I__5634\ : Odrv4
    port map (
            O => \N__31382\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__5633\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31375\
        );

    \I__5632\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31372\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31369\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__31372\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__5629\ : Odrv12
    port map (
            O => \N__31369\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__5628\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31361\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__31361\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__5626\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31354\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31351\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__31354\,
            I => \N__31348\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__31351\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__5622\ : Odrv12
    port map (
            O => \N__31348\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31343\,
            I => \N__31340\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__31340\,
            I => \N__31337\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__31337\,
            I => \N__31334\
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__31334\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__31331\,
            I => \N__31328\
        );

    \I__5616\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31325\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__31325\,
            I => \N__31322\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__31322\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__5613\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31315\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31312\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__31315\,
            I => \N__31309\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__31312\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5609\ : Odrv12
    port map (
            O => \N__31309\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__5607\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31298\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31298\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__5605\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31291\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31288\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31285\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__31288\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5601\ : Odrv12
    port map (
            O => \N__31285\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5600\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31277\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31274\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__31274\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__5597\ : CascadeMux
    port map (
            O => \N__31271\,
            I => \N__31268\
        );

    \I__5596\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31265\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__31265\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__5594\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31259\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__31259\,
            I => \N__31256\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__31256\,
            I => \N__31253\
        );

    \I__5591\ : Odrv4
    port map (
            O => \N__31253\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__31250\,
            I => \N__31247\
        );

    \I__5589\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31244\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__31244\,
            I => \N__31241\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__31241\,
            I => \N__31238\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__31238\,
            I => \N__31235\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__31235\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__5584\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31229\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__31229\,
            I => \N__31226\
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__31226\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__5580\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31217\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31214\
        );

    \I__5578\ : Span4Mux_v
    port map (
            O => \N__31214\,
            I => \N__31211\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__31211\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31205\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__31205\,
            I => \N__31202\
        );

    \I__5574\ : Odrv12
    port map (
            O => \N__31202\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__5573\ : CascadeMux
    port map (
            O => \N__31199\,
            I => \N__31196\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31193\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__5570\ : Odrv12
    port map (
            O => \N__31190\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31183\
        );

    \I__5568\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31180\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31177\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__31180\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__5565\ : Odrv12
    port map (
            O => \N__31177\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__5564\ : InMux
    port map (
            O => \N__31172\,
            I => \N__31169\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__31169\,
            I => \N__31166\
        );

    \I__5562\ : Span4Mux_v
    port map (
            O => \N__31166\,
            I => \N__31163\
        );

    \I__5561\ : Span4Mux_v
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__31160\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__5559\ : CascadeMux
    port map (
            O => \N__31157\,
            I => \N__31154\
        );

    \I__5558\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31151\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__31151\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31144\
        );

    \I__5555\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31141\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__31144\,
            I => \N__31138\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__31141\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__5552\ : Odrv12
    port map (
            O => \N__31138\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__31130\,
            I => \N__31127\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__31127\,
            I => \N__31124\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__31124\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__5547\ : CascadeMux
    port map (
            O => \N__31121\,
            I => \N__31118\
        );

    \I__5546\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31115\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__31115\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__5544\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31109\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__31109\,
            I => \N__31106\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__31106\,
            I => \N__31103\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__31103\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__5540\ : InMux
    port map (
            O => \N__31100\,
            I => \N__31097\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__31097\,
            I => \N__31093\
        );

    \I__5538\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__31090\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__31087\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__5533\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31076\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__31076\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__5531\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31070\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__31070\,
            I => \N__31067\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__31067\,
            I => \N__31064\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__31064\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__5527\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31058\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__31058\,
            I => \N__31054\
        );

    \I__5525\ : InMux
    port map (
            O => \N__31057\,
            I => \N__31051\
        );

    \I__5524\ : Span4Mux_v
    port map (
            O => \N__31054\,
            I => \N__31048\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__31051\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__5522\ : Odrv4
    port map (
            O => \N__31048\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__5520\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31037\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__31037\,
            I => \N__31034\
        );

    \I__5518\ : Odrv12
    port map (
            O => \N__31034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__5517\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31028\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__31025\,
            I => \N__31022\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__31022\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__5513\ : InMux
    port map (
            O => \N__31019\,
            I => \N__31015\
        );

    \I__5512\ : InMux
    port map (
            O => \N__31018\,
            I => \N__31012\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__31015\,
            I => \N__31009\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__31012\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__5509\ : Odrv12
    port map (
            O => \N__31009\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__5507\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30998\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__30998\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30991\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30988\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30991\,
            I => \N__30985\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__30988\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__5501\ : Odrv12
    port map (
            O => \N__30985\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__5500\ : CascadeMux
    port map (
            O => \N__30980\,
            I => \N__30977\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30974\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__30974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__30965\,
            I => \N__30962\
        );

    \I__5494\ : Span4Mux_v
    port map (
            O => \N__30962\,
            I => \N__30959\
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__30959\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30956\,
            I => \N__30952\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30949\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30952\,
            I => \N__30946\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30949\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__5488\ : Odrv12
    port map (
            O => \N__30946\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__5486\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30935\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__30935\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30925\
        );

    \I__5483\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30925\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30922\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30919\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30922\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__30919\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30914\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__5477\ : CascadeMux
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__5476\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30898\
        );

    \I__5475\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30898\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30898\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30895\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30898\,
            I => \N__30892\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30895\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__30892\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30887\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30884\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30871\
        );

    \I__5466\ : InMux
    port map (
            O => \N__30880\,
            I => \N__30871\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30871\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30868\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30871\,
            I => \N__30865\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30868\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__30865\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30857\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30857\,
            I => \N__30853\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30850\
        );

    \I__5457\ : Odrv12
    port map (
            O => \N__30853\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30850\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30842\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__30842\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__5453\ : CascadeMux
    port map (
            O => \N__30839\,
            I => \N__30836\
        );

    \I__5452\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30832\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__30835\,
            I => \N__30829\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30826\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30822\
        );

    \I__5448\ : Span4Mux_h
    port map (
            O => \N__30826\,
            I => \N__30819\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30816\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__30822\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__30819\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30816\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__5443\ : CascadeMux
    port map (
            O => \N__30809\,
            I => \N__30806\
        );

    \I__5442\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30803\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30803\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__5440\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__30797\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30790\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30787\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__30790\,
            I => \N__30784\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__30787\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__5434\ : Odrv12
    port map (
            O => \N__30784\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__30779\,
            I => \N__30776\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30776\,
            I => \N__30773\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30773\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__5430\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30767\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__30767\,
            I => \N__30763\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30760\
        );

    \I__5427\ : Span4Mux_v
    port map (
            O => \N__30763\,
            I => \N__30757\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__30760\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__30757\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30749\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__30749\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__5422\ : CascadeMux
    port map (
            O => \N__30746\,
            I => \N__30743\
        );

    \I__5421\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30740\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30740\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__30737\,
            I => \N__30734\
        );

    \I__5418\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30731\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30731\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30724\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30721\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__30724\,
            I => \N__30718\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__30721\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__5412\ : Odrv12
    port map (
            O => \N__30718\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30710\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30710\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__30707\,
            I => \N__30703\
        );

    \I__5408\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30699\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30694\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30694\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__30699\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30694\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5403\ : InMux
    port map (
            O => \N__30689\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__5401\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30677\
        );

    \I__5400\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30677\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__30677\,
            I => \N__30673\
        );

    \I__5398\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30670\
        );

    \I__5397\ : Span4Mux_h
    port map (
            O => \N__30673\,
            I => \N__30667\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__30670\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__30667\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30662\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__5393\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30652\
        );

    \I__5392\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30652\
        );

    \I__5391\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30649\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30646\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__30649\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5388\ : Odrv12
    port map (
            O => \N__30646\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5387\ : InMux
    port map (
            O => \N__30641\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__5386\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30631\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30631\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30628\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30631\,
            I => \N__30625\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__30628\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__30625\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5380\ : InMux
    port map (
            O => \N__30620\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30617\,
            I => \N__30612\
        );

    \I__5378\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30609\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30606\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__30612\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__30609\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__30606\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5373\ : InMux
    port map (
            O => \N__30599\,
            I => \bfn_11_12_0_\
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__5371\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30589\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__30592\,
            I => \N__30585\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30589\,
            I => \N__30582\
        );

    \I__5368\ : InMux
    port map (
            O => \N__30588\,
            I => \N__30579\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30576\
        );

    \I__5366\ : Span4Mux_h
    port map (
            O => \N__30582\,
            I => \N__30573\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__30579\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__30576\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__30573\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30566\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30559\
        );

    \I__5360\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30555\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30552\
        );

    \I__5358\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30549\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__30555\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__30552\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__30549\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5354\ : InMux
    port map (
            O => \N__30542\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__30539\,
            I => \N__30535\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30529\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30526\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30523\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__30526\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__30523\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30518\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30515\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30512\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30509\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30506\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__5341\ : InMux
    port map (
            O => \N__30503\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__5340\ : InMux
    port map (
            O => \N__30500\,
            I => \bfn_11_11_0_\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__30497\,
            I => \N__30493\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30496\,
            I => \N__30489\
        );

    \I__5337\ : InMux
    port map (
            O => \N__30493\,
            I => \N__30484\
        );

    \I__5336\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30484\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__30489\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__30484\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30479\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__5332\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30471\
        );

    \I__5331\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30466\
        );

    \I__5330\ : InMux
    port map (
            O => \N__30474\,
            I => \N__30466\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__30471\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__30466\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5327\ : InMux
    port map (
            O => \N__30461\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__5326\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30453\
        );

    \I__5325\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30448\
        );

    \I__5324\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30448\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__30453\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__30448\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5321\ : InMux
    port map (
            O => \N__30443\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__30440\,
            I => \N__30437\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30434\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30434\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\
        );

    \I__5317\ : InMux
    port map (
            O => \N__30431\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__5316\ : InMux
    port map (
            O => \N__30428\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__5315\ : InMux
    port map (
            O => \N__30425\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__5314\ : InMux
    port map (
            O => \N__30422\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30419\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30416\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30413\,
            I => \bfn_11_10_0_\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30410\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__5309\ : InMux
    port map (
            O => \N__30407\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30400\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30396\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__30400\,
            I => \N__30393\
        );

    \I__5305\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30390\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__30396\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__5303\ : Odrv12
    port map (
            O => \N__30393\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__30390\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__5301\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30379\
        );

    \I__5300\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30376\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__30379\,
            I => \N__30372\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__30376\,
            I => \N__30369\
        );

    \I__5297\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30365\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__30372\,
            I => \N__30360\
        );

    \I__5295\ : Span4Mux_h
    port map (
            O => \N__30369\,
            I => \N__30360\
        );

    \I__5294\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30357\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30365\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__30360\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__30357\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__30344\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df30\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__30341\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__5286\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30332\
        );

    \I__5285\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30332\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__30332\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__30329\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30323\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30323\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__5280\ : InMux
    port map (
            O => \N__30320\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__30317\,
            I => \N__30313\
        );

    \I__5278\ : CascadeMux
    port map (
            O => \N__30316\,
            I => \N__30309\
        );

    \I__5277\ : InMux
    port map (
            O => \N__30313\,
            I => \N__30302\
        );

    \I__5276\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30302\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30302\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__30302\,
            I => \N__30299\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__30299\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30293\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30290\
        );

    \I__5270\ : Span4Mux_h
    port map (
            O => \N__30290\,
            I => \N__30287\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__30287\,
            I => il_min_comp1_c
        );

    \I__5268\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__30281\,
            I => \il_max_comp1_D1\
        );

    \I__5266\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30275\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30270\
        );

    \I__5264\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30267\
        );

    \I__5263\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30264\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__30270\,
            I => \N__30260\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30257\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30254\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30263\,
            I => \N__30251\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__30260\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__30257\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__30254\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__30251\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5254\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30239\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__30239\,
            I => \N__30235\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30231\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__30235\,
            I => \N__30228\
        );

    \I__5250\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30225\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__30231\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__30228\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__30225\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__5246\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__30215\,
            I => \N__30212\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__30212\,
            I => \N__30208\
        );

    \I__5243\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30205\
        );

    \I__5242\ : Odrv4
    port map (
            O => \N__30208\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__30205\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__30200\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\
        );

    \I__5239\ : CascadeMux
    port map (
            O => \N__30197\,
            I => \N__30192\
        );

    \I__5238\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30187\
        );

    \I__5237\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30187\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30184\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__30187\,
            I => \N__30181\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__30184\,
            I => \N__30177\
        );

    \I__5233\ : Span4Mux_v
    port map (
            O => \N__30181\,
            I => \N__30174\
        );

    \I__5232\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30171\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__30177\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__30174\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__30171\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__30164\,
            I => \N__30161\
        );

    \I__5227\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30155\
        );

    \I__5226\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30155\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__30155\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30148\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30144\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__30148\,
            I => \N__30141\
        );

    \I__5221\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30138\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__30144\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__5219\ : Odrv12
    port map (
            O => \N__30141\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__30138\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__5217\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30127\
        );

    \I__5216\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30123\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30120\
        );

    \I__5214\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30117\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30114\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__30120\,
            I => \N__30108\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__30117\,
            I => \N__30108\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__30114\,
            I => \N__30105\
        );

    \I__5209\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30102\
        );

    \I__5208\ : Odrv4
    port map (
            O => \N__30108\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__30105\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__30102\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__5205\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30091\
        );

    \I__5204\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30086\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30083\
        );

    \I__5202\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30080\
        );

    \I__5201\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30077\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__30086\,
            I => \N__30073\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__30083\,
            I => \N__30070\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__30080\,
            I => \N__30065\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30065\
        );

    \I__5196\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30062\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__30073\,
            I => \N__30059\
        );

    \I__5194\ : Span4Mux_v
    port map (
            O => \N__30070\,
            I => \N__30054\
        );

    \I__5193\ : Span4Mux_h
    port map (
            O => \N__30065\,
            I => \N__30054\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__30062\,
            I => \N__30051\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__30059\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__30054\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__30051\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5188\ : InMux
    port map (
            O => \N__30044\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__30041\,
            I => \N__30038\
        );

    \I__5186\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__30029\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\
        );

    \I__5182\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30021\
        );

    \I__5181\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30018\
        );

    \I__5180\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30015\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__30021\,
            I => \N__30012\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__30018\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__30015\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__30012\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__30005\,
            I => \N__30001\
        );

    \I__5174\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29997\
        );

    \I__5173\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29994\
        );

    \I__5172\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29991\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__29997\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__29994\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29991\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__5168\ : CascadeMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29978\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__29978\,
            I => \N__29973\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29970\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29967\
        );

    \I__5163\ : Span4Mux_h
    port map (
            O => \N__29973\,
            I => \N__29962\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29957\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29967\,
            I => \N__29957\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29952\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29952\
        );

    \I__5158\ : Odrv4
    port map (
            O => \N__29962\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5157\ : Odrv12
    port map (
            O => \N__29957\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__29952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29939\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__29936\,
            I => \N__29932\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29928\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29925\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29922\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__29928\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__29925\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__29922\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__29915\,
            I => \N__29911\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29905\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29902\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29899\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29896\
        );

    \I__5140\ : InMux
    port map (
            O => \N__29908\,
            I => \N__29893\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__29905\,
            I => \N__29890\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__29902\,
            I => \N__29885\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29899\,
            I => \N__29885\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29896\,
            I => \N__29880\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29893\,
            I => \N__29880\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__29890\,
            I => \N__29875\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__29885\,
            I => \N__29875\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__29880\,
            I => \N__29872\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__29875\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__29872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__29867\,
            I => \N__29864\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29864\,
            I => \N__29861\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__29861\,
            I => \N__29858\
        );

    \I__5126\ : Span4Mux_h
    port map (
            O => \N__29858\,
            I => \N__29855\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__29855\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29846\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__29843\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__29840\,
            I => \N__29836\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29831\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29828\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__29835\,
            I => \N__29825\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__29834\,
            I => \N__29821\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29831\,
            I => \N__29818\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29815\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29812\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29809\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29806\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__29818\,
            I => \N__29801\
        );

    \I__5109\ : Span4Mux_v
    port map (
            O => \N__29815\,
            I => \N__29801\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__29812\,
            I => \N__29798\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29809\,
            I => \N__29795\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29792\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__29801\,
            I => \N__29789\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__29798\,
            I => \N__29784\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__29795\,
            I => \N__29784\
        );

    \I__5102\ : Odrv12
    port map (
            O => \N__29792\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__29789\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__29784\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5099\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__5097\ : Odrv12
    port map (
            O => \N__29771\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__5096\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29763\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29760\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29757\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__29763\,
            I => \N__29752\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29760\,
            I => \N__29749\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__29757\,
            I => \N__29746\
        );

    \I__5090\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29743\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29755\,
            I => \N__29740\
        );

    \I__5088\ : Span4Mux_v
    port map (
            O => \N__29752\,
            I => \N__29737\
        );

    \I__5087\ : Span4Mux_h
    port map (
            O => \N__29749\,
            I => \N__29734\
        );

    \I__5086\ : Span4Mux_v
    port map (
            O => \N__29746\,
            I => \N__29729\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__29743\,
            I => \N__29729\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__29740\,
            I => \N__29726\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__29737\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__29734\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__29729\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5080\ : Odrv12
    port map (
            O => \N__29726\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29714\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29711\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__29711\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__29708\,
            I => \N__29705\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29702\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__29702\,
            I => \N__29699\
        );

    \I__5073\ : Odrv12
    port map (
            O => \N__29699\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\
        );

    \I__5072\ : InMux
    port map (
            O => \N__29696\,
            I => \N__29693\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29693\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__5070\ : InMux
    port map (
            O => \N__29690\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29684\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__29684\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__5067\ : InMux
    port map (
            O => \N__29681\,
            I => \bfn_10_17_0_\
        );

    \I__5066\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29675\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__29675\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29672\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__5063\ : InMux
    port map (
            O => \N__29669\,
            I => \N__29666\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29666\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29663\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__5060\ : InMux
    port map (
            O => \N__29660\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__29654\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__5057\ : InMux
    port map (
            O => \N__29651\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__5056\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29645\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__5054\ : InMux
    port map (
            O => \N__29642\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__5053\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29636\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__29636\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__5051\ : InMux
    port map (
            O => \N__29633\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__5050\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29627\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__29627\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29624\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29618\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29618\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__5045\ : InMux
    port map (
            O => \N__29615\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__5044\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29609\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__29609\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29606\,
            I => \bfn_10_16_0_\
        );

    \I__5041\ : InMux
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__29600\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__5039\ : InMux
    port map (
            O => \N__29597\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29594\,
            I => \N__29591\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__29591\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__5036\ : InMux
    port map (
            O => \N__29588\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__5035\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__29582\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29579\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__29576\,
            I => \N__29573\
        );

    \I__5031\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29570\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__29567\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29564\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29558\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29558\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__5025\ : InMux
    port map (
            O => \N__29555\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__5024\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__29549\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29546\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29543\,
            I => \N__29540\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__29540\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__5019\ : InMux
    port map (
            O => \N__29537\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__5018\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29531\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__29531\,
            I => \N__29528\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__29528\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29525\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__5013\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__29516\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29513\,
            I => \bfn_10_15_0_\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29507\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__29507\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29504\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__5007\ : InMux
    port map (
            O => \N__29501\,
            I => \N__29498\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__29498\,
            I => \N__29495\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__29495\,
            I => \N__29492\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__29492\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__5003\ : InMux
    port map (
            O => \N__29489\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__5002\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29483\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__29483\,
            I => \N__29480\
        );

    \I__5000\ : Span4Mux_h
    port map (
            O => \N__29480\,
            I => \N__29477\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__29477\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__4998\ : InMux
    port map (
            O => \N__29474\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29468\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29468\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__4995\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29462\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__29462\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_12\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29459\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29453\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__29453\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_13\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29450\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__4989\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29440\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29440\
        );

    \I__4987\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29437\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29428\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__29434\,
            I => \N__29428\
        );

    \I__4983\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29425\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__29428\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__29425\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29420\,
            I => \N__29417\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29417\,
            I => \N__29413\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29410\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__29413\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__29410\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__4975\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29401\
        );

    \I__4974\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29398\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__29401\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__29398\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29389\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29386\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29389\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__29386\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29378\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29372\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__29372\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__4963\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__29366\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__4961\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29360\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__29360\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__4959\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29354\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__29354\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__4957\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29348\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__29348\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__4955\ : InMux
    port map (
            O => \N__29345\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__29342\,
            I => \N__29339\
        );

    \I__4953\ : InMux
    port map (
            O => \N__29339\,
            I => \N__29336\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__29336\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29333\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__4950\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29327\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29327\,
            I => \N__29322\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29319\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29316\
        );

    \I__4946\ : Span12Mux_h
    port map (
            O => \N__29322\,
            I => \N__29313\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__29319\,
            I => \N__29310\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29316\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4943\ : Odrv12
    port map (
            O => \N__29313\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__29310\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4941\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29300\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__29297\,
            I => \N__29293\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29290\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__29293\,
            I => \N__29285\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__29290\,
            I => \N__29282\
        );

    \I__4935\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29277\
        );

    \I__4934\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29277\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__29285\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4932\ : Odrv4
    port map (
            O => \N__29282\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__29277\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4930\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29267\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__29267\,
            I => \N__29262\
        );

    \I__4928\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29259\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29256\
        );

    \I__4926\ : Span12Mux_v
    port map (
            O => \N__29262\,
            I => \N__29253\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__29259\,
            I => \N__29250\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__29256\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4923\ : Odrv12
    port map (
            O => \N__29253\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__29250\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29240\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__29240\,
            I => \N__29237\
        );

    \I__4919\ : Span4Mux_v
    port map (
            O => \N__29237\,
            I => \N__29231\
        );

    \I__4918\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29228\
        );

    \I__4917\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29223\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29223\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__29231\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__29228\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__29223\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4912\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29213\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__29213\,
            I => \N__29210\
        );

    \I__4910\ : Span4Mux_h
    port map (
            O => \N__29210\,
            I => \N__29206\
        );

    \I__4909\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29202\
        );

    \I__4908\ : Span4Mux_v
    port map (
            O => \N__29206\,
            I => \N__29199\
        );

    \I__4907\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29196\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__29202\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__29199\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__29196\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4903\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29185\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29181\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29178\
        );

    \I__4900\ : CascadeMux
    port map (
            O => \N__29184\,
            I => \N__29174\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29181\,
            I => \N__29171\
        );

    \I__4898\ : Span4Mux_v
    port map (
            O => \N__29178\,
            I => \N__29168\
        );

    \I__4897\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29163\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29163\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__29171\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__29168\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__29163\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4892\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29149\
        );

    \I__4890\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29146\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__29149\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__29146\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4887\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29136\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29131\
        );

    \I__4885\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29131\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29128\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__29131\,
            I => \N__29125\
        );

    \I__4882\ : Span4Mux_h
    port map (
            O => \N__29128\,
            I => \N__29121\
        );

    \I__4881\ : Span4Mux_v
    port map (
            O => \N__29125\,
            I => \N__29118\
        );

    \I__4880\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29115\
        );

    \I__4879\ : Odrv4
    port map (
            O => \N__29121\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__29118\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__29115\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__29108\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__29105\,
            I => \N__29102\
        );

    \I__4874\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29096\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29096\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__29096\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__29090\,
            I => \N__29087\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__29087\,
            I => \N__29083\
        );

    \I__4868\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29080\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__29083\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__29080\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4865\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29068\
        );

    \I__4864\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29068\
        );

    \I__4863\ : InMux
    port map (
            O => \N__29073\,
            I => \N__29064\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29061\
        );

    \I__4861\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29058\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__29064\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__29061\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__29058\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__29051\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__29048\,
            I => \N__29045\
        );

    \I__4855\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29041\
        );

    \I__4854\ : InMux
    port map (
            O => \N__29044\,
            I => \N__29038\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__29041\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__29038\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__4851\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__29030\,
            I => \N__29027\
        );

    \I__4849\ : Span4Mux_v
    port map (
            O => \N__29027\,
            I => \N__29023\
        );

    \I__4848\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29020\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__29023\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__29020\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__29015\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\
        );

    \I__4844\ : InMux
    port map (
            O => \N__29012\,
            I => \N__29009\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__29006\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__29006\,
            I => \N__29000\
        );

    \I__4841\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28995\
        );

    \I__4840\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28995\
        );

    \I__4839\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28992\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__29000\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28995\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__28992\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28976\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28976\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__28976\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28970\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__28970\,
            I => \N__28967\
        );

    \I__4829\ : Span4Mux_h
    port map (
            O => \N__28967\,
            I => \N__28963\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28960\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__28963\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__28960\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__28955\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28949\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__28949\,
            I => \N__28944\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28939\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28939\
        );

    \I__4820\ : Span4Mux_h
    port map (
            O => \N__28944\,
            I => \N__28933\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__28939\,
            I => \N__28933\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28930\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__28933\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__28930\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28919\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28919\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__28919\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28913\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28910\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__28910\,
            I => \N__28906\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28903\
        );

    \I__4808\ : Odrv4
    port map (
            O => \N__28906\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__28903\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__28898\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28890\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28885\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28885\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28881\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28885\,
            I => \N__28878\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28875\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__28881\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__28878\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__28875\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28862\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28862\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__28862\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__28853\,
            I => \N__28848\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28845\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28842\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__28848\,
            I => \N__28839\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28845\,
            I => \N__28836\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__28842\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28839\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__28836\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4783\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28826\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__28823\,
            I => \N__28819\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28816\
        );

    \I__4779\ : Span4Mux_v
    port map (
            O => \N__28819\,
            I => \N__28811\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28808\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28803\
        );

    \I__4776\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28803\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__28811\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__28808\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__28803\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__28796\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28787\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28784\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28779\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28779\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28787\,
            I => \N__28776\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28784\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__28779\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__28776\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28765\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__28768\,
            I => \N__28762\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28765\,
            I => \N__28759\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28756\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__28759\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__28756\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__28751\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28745\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28745\,
            I => \N__28739\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28736\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28731\
        );

    \I__4752\ : InMux
    port map (
            O => \N__28742\,
            I => \N__28731\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__28739\,
            I => \N__28728\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__28736\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__28731\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__28728\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__28721\,
            I => \N__28716\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__28720\,
            I => \N__28713\
        );

    \I__4745\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28706\
        );

    \I__4744\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28706\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28706\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__28706\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28703\,
            I => \N__28694\
        );

    \I__4740\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28694\
        );

    \I__4739\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28694\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__28694\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28688\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__28688\,
            I => \N__28684\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28681\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__28684\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__28681\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__4732\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28670\
        );

    \I__4731\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28665\
        );

    \I__4730\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28665\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28662\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__28670\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__28665\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28662\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__4725\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28651\
        );

    \I__4724\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28646\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28643\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28638\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28638\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__28646\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__28643\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__28638\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28626\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28623\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28629\,
            I => \N__28620\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28626\,
            I => \N__28617\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28614\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__28620\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__28617\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__4710\ : Odrv12
    port map (
            O => \N__28614\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28599\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28599\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__28605\,
            I => \N__28596\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28593\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28590\
        );

    \I__4704\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28587\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__28593\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__28590\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28587\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28577\,
            I => \N__28574\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__28574\,
            I => \N__28570\
        );

    \I__4697\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28567\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__28570\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__28567\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28559\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28559\,
            I => \N__28554\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28551\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__28557\,
            I => \N__28548\
        );

    \I__4690\ : Span4Mux_v
    port map (
            O => \N__28554\,
            I => \N__28542\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28542\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28539\
        );

    \I__4687\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28536\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__28542\,
            I => \N__28533\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28530\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__28536\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__28533\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__28530\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__28523\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28517\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__28514\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__4677\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28508\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__28508\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__28502\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__4673\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28496\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__28496\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28490\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28486\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28483\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__28486\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__28483\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__28478\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__4663\ : Odrv12
    port map (
            O => \N__28469\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__28466\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__4661\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28459\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28456\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28451\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28456\,
            I => \N__28448\
        );

    \I__4657\ : InMux
    port map (
            O => \N__28455\,
            I => \N__28443\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28454\,
            I => \N__28443\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__28451\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__28448\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__28443\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__28436\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28426\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28423\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__28426\,
            I => \N__28417\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28417\
        );

    \I__4646\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28414\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__28417\,
            I => \N__28411\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__28414\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__28411\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4642\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28403\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__4640\ : Span4Mux_v
    port map (
            O => \N__28400\,
            I => \N__28396\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28399\,
            I => \N__28393\
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__28396\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__28393\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__28388\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28382\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__28382\,
            I => \N__28376\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28373\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28368\
        );

    \I__4631\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28368\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__28376\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28373\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__28368\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4627\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28358\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28355\,
            I => \N__28352\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__28352\,
            I => \N__28348\
        );

    \I__4623\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__28348\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__28345\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__28340\,
            I => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28331\
        );

    \I__4618\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28324\
        );

    \I__4617\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28324\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28324\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__28331\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__28324\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__28319\,
            I => \N__28316\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28310\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__28310\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__4609\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28304\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__28304\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28298\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28294\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__28297\,
            I => \N__28289\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__28294\,
            I => \N__28286\
        );

    \I__4603\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28283\
        );

    \I__4602\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28280\
        );

    \I__4601\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28277\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__28286\,
            I => \N__28272\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__28283\,
            I => \N__28272\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__28280\,
            I => \N__28269\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__28277\,
            I => \N__28264\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__28272\,
            I => \N__28264\
        );

    \I__4595\ : Span4Mux_h
    port map (
            O => \N__28269\,
            I => \N__28261\
        );

    \I__4594\ : Span4Mux_h
    port map (
            O => \N__28264\,
            I => \N__28258\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__28261\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__28258\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__28253\,
            I => \N__28250\
        );

    \I__4590\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28247\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28247\,
            I => \N__28244\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__28244\,
            I => \N__28241\
        );

    \I__4587\ : Span4Mux_h
    port map (
            O => \N__28241\,
            I => \N__28238\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__28238\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__28235\,
            I => \N__28230\
        );

    \I__4584\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28226\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28223\
        );

    \I__4582\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28220\
        );

    \I__4581\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28217\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__28226\,
            I => \N__28214\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__28223\,
            I => \N__28209\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28209\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28206\
        );

    \I__4576\ : Span4Mux_h
    port map (
            O => \N__28214\,
            I => \N__28200\
        );

    \I__4575\ : Span4Mux_h
    port map (
            O => \N__28209\,
            I => \N__28200\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__28206\,
            I => \N__28197\
        );

    \I__4573\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28194\
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__28200\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__28197\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__28194\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4569\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28183\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__28186\,
            I => \N__28180\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28176\
        );

    \I__4566\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28171\
        );

    \I__4565\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28171\
        );

    \I__4564\ : Span4Mux_h
    port map (
            O => \N__28176\,
            I => \N__28166\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28166\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__28166\,
            I => \N__28163\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__28163\,
            I => \N__28160\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__28160\,
            I => \N__28157\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__28157\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4558\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28147\
        );

    \I__4556\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28144\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__28147\,
            I => \N__28139\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__28144\,
            I => \N__28139\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__28139\,
            I => \N__28136\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__28136\,
            I => \N__28131\
        );

    \I__4551\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28126\
        );

    \I__4550\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28126\
        );

    \I__4549\ : Span4Mux_v
    port map (
            O => \N__28131\,
            I => \N__28123\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__28126\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__28123\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4546\ : ClkMux
    port map (
            O => \N__28118\,
            I => \N__28115\
        );

    \I__4545\ : GlobalMux
    port map (
            O => \N__28115\,
            I => \N__28112\
        );

    \I__4544\ : gio2CtrlBuf
    port map (
            O => \N__28112\,
            I => delay_tr_input_c_g
        );

    \I__4543\ : IoInMux
    port map (
            O => \N__28109\,
            I => \N__28106\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__28106\,
            I => \N__28103\
        );

    \I__4541\ : Odrv12
    port map (
            O => \N__28103\,
            I => s3_phy_c
        );

    \I__4540\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28097\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__4538\ : Glb2LocalMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__4537\ : GlobalMux
    port map (
            O => \N__28091\,
            I => clk_12mhz
        );

    \I__4536\ : IoInMux
    port map (
            O => \N__28088\,
            I => \N__28085\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__28085\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__4534\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__4532\ : Span4Mux_h
    port map (
            O => \N__28076\,
            I => \N__28073\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__28073\,
            I => il_max_comp1_c
        );

    \I__4530\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__28067\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4527\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28057\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__28060\,
            I => \N__28054\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28049\
        );

    \I__4524\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28044\
        );

    \I__4523\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28044\
        );

    \I__4522\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28040\
        );

    \I__4521\ : Span4Mux_v
    port map (
            O => \N__28049\,
            I => \N__28035\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__28044\,
            I => \N__28035\
        );

    \I__4519\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28032\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__28040\,
            I => \N__28027\
        );

    \I__4517\ : Span4Mux_h
    port map (
            O => \N__28035\,
            I => \N__28027\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__28032\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__28027\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__28022\,
            I => \N__28019\
        );

    \I__4513\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__28016\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\
        );

    \I__4511\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28008\
        );

    \I__4510\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28005\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__28011\,
            I => \N__28001\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__27998\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__28005\,
            I => \N__27995\
        );

    \I__4506\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27991\
        );

    \I__4505\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27988\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__27998\,
            I => \N__27983\
        );

    \I__4503\ : Span4Mux_v
    port map (
            O => \N__27995\,
            I => \N__27983\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27980\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__27991\,
            I => \N__27975\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27975\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__27983\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__27980\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4497\ : Odrv12
    port map (
            O => \N__27975\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27962\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__4491\ : Odrv4
    port map (
            O => \N__27953\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__27950\,
            I => \N__27946\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27943\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27940\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27943\,
            I => \N__27935\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27932\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27926\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27926\
        );

    \I__4483\ : Span4Mux_h
    port map (
            O => \N__27935\,
            I => \N__27921\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__27932\,
            I => \N__27921\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27918\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27915\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__27921\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27918\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__27915\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__27908\,
            I => \N__27905\
        );

    \I__4475\ : InMux
    port map (
            O => \N__27905\,
            I => \N__27902\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__27902\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__27893\,
            I => \N__27890\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__27890\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__27887\,
            I => \N__27884\
        );

    \I__4468\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27881\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27881\,
            I => \N__27878\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__27878\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\
        );

    \I__4465\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27872\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27869\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__27869\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__27866\,
            I => \N__27863\
        );

    \I__4461\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27858\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27855\
        );

    \I__4459\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27851\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27846\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27846\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27843\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27851\,
            I => \N__27838\
        );

    \I__4454\ : Span4Mux_h
    port map (
            O => \N__27846\,
            I => \N__27838\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27843\,
            I => \N__27832\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__27838\,
            I => \N__27832\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27829\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__27832\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27829\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27821\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27821\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27814\
        );

    \I__4445\ : CascadeMux
    port map (
            O => \N__27817\,
            I => \N__27810\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27805\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27802\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27799\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27796\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27793\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__27805\,
            I => \N__27790\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27783\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27783\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27783\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27780\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__27790\,
            I => \N__27775\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__27783\,
            I => \N__27775\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__27780\,
            I => \N__27772\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__27775\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__27772\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27764\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__27761\,
            I => \N__27758\
        );

    \I__4426\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27752\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__27752\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__27749\,
            I => \N__27745\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27740\
        );

    \I__4421\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27737\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27734\
        );

    \I__4419\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27730\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27740\,
            I => \N__27727\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__27737\,
            I => \N__27722\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27722\
        );

    \I__4415\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27719\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__27730\,
            I => \N__27716\
        );

    \I__4413\ : Span12Mux_h
    port map (
            O => \N__27727\,
            I => \N__27709\
        );

    \I__4412\ : Span12Mux_s7_h
    port map (
            O => \N__27722\,
            I => \N__27709\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27719\,
            I => \N__27709\
        );

    \I__4410\ : Odrv12
    port map (
            O => \N__27716\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4409\ : Odrv12
    port map (
            O => \N__27709\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27698\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27689\
        );

    \I__4404\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27686\
        );

    \I__4403\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27680\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27680\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__27689\,
            I => \N__27677\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27674\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27671\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27680\,
            I => \N__27668\
        );

    \I__4397\ : Span4Mux_h
    port map (
            O => \N__27677\,
            I => \N__27665\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__27674\,
            I => \N__27658\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__27671\,
            I => \N__27658\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__27668\,
            I => \N__27658\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__27665\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__27658\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__27653\,
            I => \N__27650\
        );

    \I__4390\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27647\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27641\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__27641\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__27638\,
            I => \N__27635\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27631\
        );

    \I__4384\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27625\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__27631\,
            I => \N__27622\
        );

    \I__4382\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27617\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27617\
        );

    \I__4380\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27614\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__27625\,
            I => \N__27611\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__27622\,
            I => \N__27608\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__27617\,
            I => \N__27605\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__27614\,
            I => \N__27602\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__27611\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__27608\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__27605\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4372\ : Odrv12
    port map (
            O => \N__27602\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__27593\,
            I => \N__27590\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27587\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__27587\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27581\,
            I => \N__27578\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__27578\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\
        );

    \I__4365\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27571\
        );

    \I__4364\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27568\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__27571\,
            I => \N__27564\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__27568\,
            I => \N__27561\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27556\
        );

    \I__4360\ : Span4Mux_h
    port map (
            O => \N__27564\,
            I => \N__27551\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__27561\,
            I => \N__27551\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27546\
        );

    \I__4357\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27546\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__27556\,
            I => \N__27543\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__27551\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27546\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__27543\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4352\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27533\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__27530\,
            I => \N__27525\
        );

    \I__4349\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27522\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27519\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27515\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27512\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27519\,
            I => \N__27509\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27506\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__27515\,
            I => \N__27503\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__27512\,
            I => \N__27500\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__27509\,
            I => \N__27496\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27493\
        );

    \I__4339\ : Span4Mux_v
    port map (
            O => \N__27503\,
            I => \N__27488\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__27500\,
            I => \N__27488\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27485\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__27496\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4335\ : Odrv12
    port map (
            O => \N__27493\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__27488\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27485\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__4331\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27470\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__27470\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27467\,
            I => \N__27464\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__27464\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__27461\,
            I => \N__27458\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27455\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__27455\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__27452\,
            I => \N__27449\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27446\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__27446\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__27443\,
            I => \N__27440\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27437\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__27437\,
            I => \N__27434\
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__27434\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \N__27427\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__27430\,
            I => \N__27424\
        );

    \I__4315\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27419\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27416\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27413\
        );

    \I__4312\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27410\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27404\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27404\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__27413\,
            I => \N__27401\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27398\
        );

    \I__4307\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27395\
        );

    \I__4306\ : Span4Mux_v
    port map (
            O => \N__27404\,
            I => \N__27388\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__27401\,
            I => \N__27388\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__27398\,
            I => \N__27388\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27383\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__27388\,
            I => \N__27383\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__27383\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__27380\,
            I => \N__27377\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27374\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__27374\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27366\
        );

    \I__4296\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27362\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__27369\,
            I => \N__27359\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__27366\,
            I => \N__27356\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27353\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27349\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27346\
        );

    \I__4290\ : Span4Mux_v
    port map (
            O => \N__27356\,
            I => \N__27341\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__27353\,
            I => \N__27341\
        );

    \I__4288\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27338\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__27349\,
            I => \N__27335\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__27346\,
            I => \N__27330\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__27341\,
            I => \N__27330\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__27338\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__27335\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__27330\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__4280\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27317\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27314\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__27314\,
            I => \N__27311\
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__27311\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__4275\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27302\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__27302\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\
        );

    \I__4273\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__27293\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__4270\ : CascadeMux
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__4269\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27284\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27284\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\
        );

    \I__4267\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27278\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__27278\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__4264\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27268\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27265\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__27268\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_14\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27265\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_14\
        );

    \I__4260\ : CascadeMux
    port map (
            O => \N__27260\,
            I => \N__27256\
        );

    \I__4259\ : InMux
    port map (
            O => \N__27259\,
            I => \N__27253\
        );

    \I__4258\ : InMux
    port map (
            O => \N__27256\,
            I => \N__27250\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__27253\,
            I => \N__27247\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__27250\,
            I => \N__27242\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__27247\,
            I => \N__27242\
        );

    \I__4254\ : Span4Mux_h
    port map (
            O => \N__27242\,
            I => \N__27237\
        );

    \I__4253\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27232\
        );

    \I__4252\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27232\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__27237\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__27232\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4249\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27224\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27224\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__27221\,
            I => \N__27218\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4244\ : Span4Mux_h
    port map (
            O => \N__27212\,
            I => \N__27209\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__27209\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \N__27203\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27197\
        );

    \I__4240\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27194\
        );

    \I__4239\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27190\
        );

    \I__4238\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27187\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__27197\,
            I => \N__27184\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__27194\,
            I => \N__27181\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27178\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__27190\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__27187\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__27184\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__27181\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__27178\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__27167\,
            I => \N__27164\
        );

    \I__4228\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27161\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__27161\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__27158\,
            I => \N__27154\
        );

    \I__4225\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27150\
        );

    \I__4224\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27146\
        );

    \I__4223\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27143\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27140\
        );

    \I__4221\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27137\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27132\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__27143\,
            I => \N__27132\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__27140\,
            I => \N__27126\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__27137\,
            I => \N__27126\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__27132\,
            I => \N__27123\
        );

    \I__4215\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27120\
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__27126\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__27123\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__27120\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__4210\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__27107\,
            I => \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\
        );

    \I__4208\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27100\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__27103\,
            I => \N__27097\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27094\
        );

    \I__4205\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27091\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__27094\,
            I => \N__27088\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27085\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__27088\,
            I => \N__27080\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__27085\,
            I => \N__27077\
        );

    \I__4200\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27072\
        );

    \I__4199\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27072\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__27080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__27077\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__27072\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__27065\,
            I => \N__27062\
        );

    \I__4194\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27059\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__27059\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__27056\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__4190\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27045\
        );

    \I__4189\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27040\
        );

    \I__4188\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27040\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__27045\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__27040\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4185\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27030\
        );

    \I__4184\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27025\
        );

    \I__4183\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27025\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27022\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__27025\,
            I => \N__27019\
        );

    \I__4180\ : Span4Mux_h
    port map (
            O => \N__27022\,
            I => \N__27016\
        );

    \I__4179\ : Span12Mux_h
    port map (
            O => \N__27019\,
            I => \N__27013\
        );

    \I__4178\ : Span4Mux_v
    port map (
            O => \N__27016\,
            I => \N__27010\
        );

    \I__4177\ : Span12Mux_v
    port map (
            O => \N__27013\,
            I => \N__27007\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__27010\,
            I => \N__27004\
        );

    \I__4175\ : Odrv12
    port map (
            O => \N__27007\,
            I => il_min_comp2_c
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__27004\,
            I => il_min_comp2_c
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__26999\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2_cascade_\
        );

    \I__4172\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__4170\ : Sp12to4
    port map (
            O => \N__26990\,
            I => \N__26984\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26979\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26979\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26976\
        );

    \I__4166\ : Odrv12
    port map (
            O => \N__26984\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26979\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__26976\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26966\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__26963\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__26960\,
            I => \N__26956\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26953\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26950\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26945\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26950\,
            I => \N__26945\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__26942\,
            I => \N__26938\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26935\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__26938\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26935\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26927\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__26924\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__26921\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0_cascade_\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26912\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__26909\,
            I => \N__26906\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__26906\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26900\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__26897\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__4138\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26891\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26887\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26884\
        );

    \I__4135\ : Odrv12
    port map (
            O => \N__26887\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26884\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__26879\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26876\,
            I => \N__26872\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26869\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26872\,
            I => \N__26866\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26861\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__26866\,
            I => \N__26858\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26853\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26853\
        );

    \I__4125\ : Span4Mux_h
    port map (
            O => \N__26861\,
            I => \N__26850\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__26858\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26853\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__26850\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__26843\,
            I => \N__26839\
        );

    \I__4120\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26834\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26834\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26834\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26828\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__26828\,
            I => \N__26823\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26820\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26817\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__26823\,
            I => \N__26814\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26811\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26817\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__26814\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4109\ : Odrv12
    port map (
            O => \N__26811\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26798\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26798\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__26798\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26792\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26792\,
            I => \N__26788\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26782\
        );

    \I__4102\ : Span4Mux_h
    port map (
            O => \N__26788\,
            I => \N__26779\
        );

    \I__4101\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26772\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26772\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26772\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26782\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__26779\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26772\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26759\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26759\,
            I => \N__26755\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26752\
        );

    \I__4091\ : Span4Mux_v
    port map (
            O => \N__26755\,
            I => \N__26749\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26752\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__26749\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__26744\,
            I => \N__26740\
        );

    \I__4087\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26737\
        );

    \I__4086\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26733\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__26737\,
            I => \N__26730\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26725\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26733\,
            I => \N__26722\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__26730\,
            I => \N__26719\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26714\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26714\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__26725\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__26722\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__26719\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__26714\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26696\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26696\
        );

    \I__4073\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26696\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26696\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26686\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26683\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__26686\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__26683\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4066\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26675\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__26675\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26672\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__26669\,
            I => \N__26666\
        );

    \I__4062\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26662\
        );

    \I__4061\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26659\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26653\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26653\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26650\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__26653\,
            I => \N__26647\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__26650\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__26647\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26642\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__26639\,
            I => \N__26635\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__26638\,
            I => \N__26632\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26629\
        );

    \I__4050\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26626\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26629\,
            I => \N__26620\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__26626\,
            I => \N__26620\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26617\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26617\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__26614\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4043\ : InMux
    port map (
            O => \N__26609\,
            I => \bfn_9_11_0_\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26598\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26595\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26592\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__26598\,
            I => \N__26587\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__26595\,
            I => \N__26587\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26592\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4035\ : Odrv12
    port map (
            O => \N__26587\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26582\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26572\
        );

    \I__4032\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26572\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26569\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__26572\,
            I => \N__26566\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__26569\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4028\ : Odrv12
    port map (
            O => \N__26566\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4027\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__4026\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26554\
        );

    \I__4025\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26551\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26548\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__26551\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__4022\ : Odrv12
    port map (
            O => \N__26548\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__4021\ : InMux
    port map (
            O => \N__26543\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26533\
        );

    \I__4018\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26530\
        );

    \I__4017\ : Span4Mux_v
    port map (
            O => \N__26533\,
            I => \N__26527\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__26530\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__26527\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__26522\,
            I => \N__26519\
        );

    \I__4013\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26514\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26511\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26508\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__26514\,
            I => \N__26503\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__26511\,
            I => \N__26503\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__26508\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4007\ : Odrv12
    port map (
            O => \N__26503\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4006\ : InMux
    port map (
            O => \N__26498\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26495\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__4004\ : CEMux
    port map (
            O => \N__26492\,
            I => \N__26487\
        );

    \I__4003\ : CEMux
    port map (
            O => \N__26491\,
            I => \N__26484\
        );

    \I__4002\ : CEMux
    port map (
            O => \N__26490\,
            I => \N__26480\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__26487\,
            I => \N__26476\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26484\,
            I => \N__26473\
        );

    \I__3999\ : CEMux
    port map (
            O => \N__26483\,
            I => \N__26470\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__26480\,
            I => \N__26467\
        );

    \I__3997\ : CEMux
    port map (
            O => \N__26479\,
            I => \N__26464\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__26476\,
            I => \N__26457\
        );

    \I__3995\ : Span4Mux_v
    port map (
            O => \N__26473\,
            I => \N__26457\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26470\,
            I => \N__26457\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__26467\,
            I => \N__26454\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__26464\,
            I => \N__26451\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__26457\,
            I => \delay_measurement_inst.delay_tr_timer.N_203_i\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__26454\,
            I => \delay_measurement_inst.delay_tr_timer.N_203_i\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__26451\,
            I => \delay_measurement_inst.delay_tr_timer.N_203_i\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26440\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26443\,
            I => \N__26437\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__26440\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26437\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26428\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26425\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__26428\,
            I => \N__26420\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__26425\,
            I => \N__26417\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26412\
        );

    \I__3979\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26412\
        );

    \I__3978\ : Span4Mux_v
    port map (
            O => \N__26420\,
            I => \N__26407\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__26417\,
            I => \N__26407\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__26412\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__26407\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__26402\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26393\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26398\,
            I => \N__26393\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26393\,
            I => \N__26389\
        );

    \I__3970\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26386\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__26389\,
            I => \N__26383\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__26386\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__26383\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26378\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__26375\,
            I => \N__26371\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__26374\,
            I => \N__26368\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26362\
        );

    \I__3962\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26362\
        );

    \I__3961\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26359\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26362\,
            I => \N__26356\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__26359\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3958\ : Odrv12
    port map (
            O => \N__26356\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3957\ : InMux
    port map (
            O => \N__26351\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__26348\,
            I => \N__26344\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__26347\,
            I => \N__26341\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26338\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26335\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26338\,
            I => \N__26329\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__26335\,
            I => \N__26329\
        );

    \I__3950\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26326\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__26329\,
            I => \N__26323\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26326\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__26323\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3946\ : InMux
    port map (
            O => \N__26318\,
            I => \bfn_9_10_0_\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__3944\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26304\
        );

    \I__3942\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26301\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26307\,
            I => \N__26298\
        );

    \I__3940\ : Sp12to4
    port map (
            O => \N__26304\,
            I => \N__26293\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__26301\,
            I => \N__26293\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__26298\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3937\ : Odrv12
    port map (
            O => \N__26293\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26288\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__3935\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26278\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26278\
        );

    \I__3933\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26275\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__26278\,
            I => \N__26272\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__26275\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3930\ : Odrv12
    port map (
            O => \N__26272\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3929\ : InMux
    port map (
            O => \N__26267\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26257\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26257\
        );

    \I__3926\ : InMux
    port map (
            O => \N__26262\,
            I => \N__26254\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26251\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__26254\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3923\ : Odrv12
    port map (
            O => \N__26251\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26246\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__26243\,
            I => \N__26239\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__26242\,
            I => \N__26236\
        );

    \I__3919\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26230\
        );

    \I__3918\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26230\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26227\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26224\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__26227\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3914\ : Odrv12
    port map (
            O => \N__26224\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3913\ : InMux
    port map (
            O => \N__26219\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__26216\,
            I => \N__26212\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \N__26209\
        );

    \I__3910\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26203\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26203\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26200\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26197\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26200\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3905\ : Odrv12
    port map (
            O => \N__26197\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3904\ : InMux
    port map (
            O => \N__26192\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3903\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26183\
        );

    \I__3902\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26183\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26179\
        );

    \I__3900\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26176\
        );

    \I__3899\ : Span4Mux_v
    port map (
            O => \N__26179\,
            I => \N__26173\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__26176\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3897\ : Odrv4
    port map (
            O => \N__26173\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3896\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26162\
        );

    \I__3895\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26162\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__26162\,
            I => \N__26158\
        );

    \I__3893\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26155\
        );

    \I__3892\ : Span4Mux_v
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__26155\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__26152\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3889\ : InMux
    port map (
            O => \N__26147\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3888\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__3887\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26138\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26134\
        );

    \I__3885\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26131\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__26134\,
            I => \N__26128\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__26131\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__26128\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3881\ : InMux
    port map (
            O => \N__26123\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__26120\,
            I => \N__26116\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__26119\,
            I => \N__26113\
        );

    \I__3878\ : InMux
    port map (
            O => \N__26116\,
            I => \N__26110\
        );

    \I__3877\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26107\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26110\,
            I => \N__26101\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26101\
        );

    \I__3874\ : InMux
    port map (
            O => \N__26106\,
            I => \N__26098\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__26101\,
            I => \N__26095\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__26098\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__26095\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3870\ : InMux
    port map (
            O => \N__26090\,
            I => \bfn_9_9_0_\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__26087\,
            I => \N__26083\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__26086\,
            I => \N__26080\
        );

    \I__3867\ : InMux
    port map (
            O => \N__26083\,
            I => \N__26076\
        );

    \I__3866\ : InMux
    port map (
            O => \N__26080\,
            I => \N__26073\
        );

    \I__3865\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26070\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26065\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__26073\,
            I => \N__26065\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__26070\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3861\ : Odrv12
    port map (
            O => \N__26065\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3860\ : InMux
    port map (
            O => \N__26060\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__3859\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26051\
        );

    \I__3858\ : InMux
    port map (
            O => \N__26056\,
            I => \N__26051\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__26051\,
            I => \N__26047\
        );

    \I__3856\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26044\
        );

    \I__3855\ : Span4Mux_v
    port map (
            O => \N__26047\,
            I => \N__26041\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__26044\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__26041\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3852\ : InMux
    port map (
            O => \N__26036\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__3850\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26026\
        );

    \I__3849\ : InMux
    port map (
            O => \N__26029\,
            I => \N__26023\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__26026\,
            I => \N__26017\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__26023\,
            I => \N__26017\
        );

    \I__3846\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26014\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__26017\,
            I => \N__26011\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__26014\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__26011\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3842\ : InMux
    port map (
            O => \N__26006\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__26003\,
            I => \N__25999\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__26002\,
            I => \N__25996\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25990\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25990\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25987\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25990\,
            I => \N__25984\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25987\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3834\ : Odrv12
    port map (
            O => \N__25984\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25979\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25969\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25969\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25966\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25969\,
            I => \N__25963\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25966\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3827\ : Odrv12
    port map (
            O => \N__25963\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25958\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25955\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25952\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__3823\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25911\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25911\
        );

    \I__3821\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25911\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25911\
        );

    \I__3819\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25902\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25902\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25902\
        );

    \I__3816\ : InMux
    port map (
            O => \N__25942\,
            I => \N__25902\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25893\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25893\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25893\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25893\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25888\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25888\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25879\
        );

    \I__3808\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25879\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25879\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25879\
        );

    \I__3805\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25870\
        );

    \I__3804\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25870\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25870\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25870\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25861\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25861\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25861\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25861\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25923\,
            I => \N__25852\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25852\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25852\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25920\,
            I => \N__25852\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25911\,
            I => \N__25845\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25845\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25893\,
            I => \N__25845\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25888\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__25879\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25870\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25861\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25852\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__25845\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3784\ : InMux
    port map (
            O => \N__25832\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__3783\ : CEMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__25826\,
            I => \N__25822\
        );

    \I__3781\ : CEMux
    port map (
            O => \N__25825\,
            I => \N__25819\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__25822\,
            I => \N__25813\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25819\,
            I => \N__25813\
        );

    \I__3778\ : CEMux
    port map (
            O => \N__25818\,
            I => \N__25810\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__25813\,
            I => \N__25806\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__25810\,
            I => \N__25803\
        );

    \I__3775\ : CEMux
    port map (
            O => \N__25809\,
            I => \N__25800\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__25806\,
            I => \N__25795\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__25803\,
            I => \N__25795\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25800\,
            I => \N__25792\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__25795\,
            I => \delay_measurement_inst.delay_tr_timer.N_204_i\
        );

    \I__3770\ : Odrv12
    port map (
            O => \N__25792\,
            I => \delay_measurement_inst.delay_tr_timer.N_204_i\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__25787\,
            I => \N__25783\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25780\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25777\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__25780\,
            I => \N__25771\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__25777\,
            I => \N__25771\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25776\,
            I => \N__25768\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__25768\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__25765\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25757\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25757\,
            I => \N__25753\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25750\
        );

    \I__3757\ : Sp12to4
    port map (
            O => \N__25753\,
            I => \N__25744\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25744\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25741\
        );

    \I__3754\ : Odrv12
    port map (
            O => \N__25744\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__25741\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25736\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25727\
        );

    \I__3750\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25727\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25723\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25720\
        );

    \I__3747\ : Span4Mux_v
    port map (
            O => \N__25723\,
            I => \N__25717\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25720\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__25717\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3744\ : InMux
    port map (
            O => \N__25712\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__25709\,
            I => \N__25705\
        );

    \I__3742\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25702\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25699\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25695\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25692\
        );

    \I__3738\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25689\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__25695\,
            I => \N__25684\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__25692\,
            I => \N__25684\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__25689\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__25684\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25679\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__25676\,
            I => \N__25672\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__25675\,
            I => \N__25669\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25663\
        );

    \I__3729\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25663\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25660\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25663\,
            I => \N__25657\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__25660\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3725\ : Odrv12
    port map (
            O => \N__25657\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25652\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__25649\,
            I => \N__25645\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__25648\,
            I => \N__25642\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25645\,
            I => \N__25636\
        );

    \I__3720\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25636\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25633\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25630\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__25633\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3716\ : Odrv12
    port map (
            O => \N__25630\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3715\ : InMux
    port map (
            O => \N__25625\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3714\ : InMux
    port map (
            O => \N__25622\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25619\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25616\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__3711\ : InMux
    port map (
            O => \N__25613\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__3710\ : InMux
    port map (
            O => \N__25610\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25607\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25604\,
            I => \bfn_9_7_0_\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25601\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__3706\ : InMux
    port map (
            O => \N__25598\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25595\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__3704\ : InMux
    port map (
            O => \N__25592\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25589\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__3702\ : InMux
    port map (
            O => \N__25586\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25583\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25580\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25577\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__3698\ : InMux
    port map (
            O => \N__25574\,
            I => \bfn_9_6_0_\
        );

    \I__3697\ : InMux
    port map (
            O => \N__25571\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25568\,
            I => \bfn_9_4_0_\
        );

    \I__3695\ : InMux
    port map (
            O => \N__25565\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__3694\ : InMux
    port map (
            O => \N__25562\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__3693\ : InMux
    port map (
            O => \N__25559\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__3692\ : InMux
    port map (
            O => \N__25556\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25553\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__3690\ : InMux
    port map (
            O => \N__25550\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25547\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__3688\ : InMux
    port map (
            O => \N__25544\,
            I => \bfn_9_5_0_\
        );

    \I__3687\ : InMux
    port map (
            O => \N__25541\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__3686\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__25535\,
            I => \N__25532\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__25532\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25529\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25526\,
            I => \bfn_8_20_0_\
        );

    \I__3681\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25520\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__25514\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__25505\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__25502\,
            I => \N__25499\
        );

    \I__3673\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25495\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25498\,
            I => \N__25492\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25488\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__25492\,
            I => \N__25484\
        );

    \I__3669\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25481\
        );

    \I__3668\ : Span4Mux_v
    port map (
            O => \N__25488\,
            I => \N__25478\
        );

    \I__3667\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25475\
        );

    \I__3666\ : Span4Mux_v
    port map (
            O => \N__25484\,
            I => \N__25472\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25481\,
            I => \N__25469\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__25478\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__25475\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__25472\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__25469\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3660\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25457\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__25457\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25448\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__25448\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3655\ : IoInMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__3653\ : Odrv12
    port map (
            O => \N__25439\,
            I => s4_phy_c
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__25436\,
            I => \N__25433\
        );

    \I__3651\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25430\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__25430\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25427\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__3648\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25421\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__25421\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25418\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__25409\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3642\ : InMux
    port map (
            O => \N__25406\,
            I => \bfn_8_19_0_\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25403\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25394\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__25394\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25391\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__3635\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__25382\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3633\ : InMux
    port map (
            O => \N__25379\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__3632\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25370\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__25370\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__3629\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25364\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__25364\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25361\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__25355\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25352\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__3623\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25346\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__25346\,
            I => \N__25343\
        );

    \I__3621\ : Odrv12
    port map (
            O => \N__25343\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25340\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__3619\ : InMux
    port map (
            O => \N__25337\,
            I => \N__25334\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__3617\ : Odrv12
    port map (
            O => \N__25331\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3616\ : InMux
    port map (
            O => \N__25328\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__3615\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__3613\ : Span12Mux_v
    port map (
            O => \N__25319\,
            I => \N__25316\
        );

    \I__3612\ : Odrv12
    port map (
            O => \N__25316\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__3611\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__25310\,
            I => \N__25307\
        );

    \I__3609\ : Odrv12
    port map (
            O => \N__25307\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3608\ : InMux
    port map (
            O => \N__25304\,
            I => \bfn_8_18_0_\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__25298\,
            I => \N__25295\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__25295\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25292\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25286\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25283\
        );

    \I__3601\ : Odrv12
    port map (
            O => \N__25283\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__25280\,
            I => \N__25277\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25274\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__25271\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25268\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__3595\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__25262\,
            I => \N__25259\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__25253\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__25247\,
            I => \N__25244\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__25244\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25241\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__25238\,
            I => \N__25235\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__25229\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25226\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__25220\,
            I => \N__25217\
        );

    \I__3579\ : Span4Mux_v
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__25214\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__3577\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__25208\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3575\ : InMux
    port map (
            O => \N__25205\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__3574\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25199\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__25196\,
            I => \N__25193\
        );

    \I__3571\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__25190\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3569\ : InMux
    port map (
            O => \N__25187\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__3568\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__25178\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__25175\,
            I => \N__25172\
        );

    \I__3564\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3562\ : Span4Mux_h
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__25163\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__3560\ : InMux
    port map (
            O => \N__25160\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25157\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25151\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__25151\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25145\,
            I => \N__25142\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__25142\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__3552\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__25133\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25130\,
            I => \bfn_8_17_0_\
        );

    \I__3549\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__25121\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__3546\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__25112\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25109\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__3542\ : InMux
    port map (
            O => \N__25106\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__3541\ : InMux
    port map (
            O => \N__25103\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__3540\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__25094\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25091\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__3536\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__3534\ : Odrv12
    port map (
            O => \N__25082\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__3533\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__25070\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3529\ : InMux
    port map (
            O => \N__25067\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__3528\ : InMux
    port map (
            O => \N__25064\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__3527\ : InMux
    port map (
            O => \N__25061\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__3526\ : InMux
    port map (
            O => \N__25058\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__3525\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__25049\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__3521\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25040\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__25034\,
            I => \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\
        );

    \I__3517\ : InMux
    port map (
            O => \N__25031\,
            I => \N__25028\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__25025\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__3514\ : InMux
    port map (
            O => \N__25022\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__25019\,
            I => \N__25015\
        );

    \I__3512\ : InMux
    port map (
            O => \N__25018\,
            I => \N__25012\
        );

    \I__3511\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__25005\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__25009\,
            I => \N__25002\
        );

    \I__3508\ : InMux
    port map (
            O => \N__25008\,
            I => \N__24999\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__25005\,
            I => \N__24994\
        );

    \I__3506\ : Span4Mux_h
    port map (
            O => \N__25002\,
            I => \N__24994\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__24999\,
            I => \N__24989\
        );

    \I__3504\ : Span4Mux_h
    port map (
            O => \N__24994\,
            I => \N__24986\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24981\
        );

    \I__3502\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24981\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__24989\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__24986\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__24981\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24971\,
            I => \N__24968\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__24968\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24959\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24959\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__24956\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24948\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24943\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24943\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__24948\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__24943\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__24938\,
            I => \N__24935\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24928\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24928\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24925\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24925\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__24922\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__24917\,
            I => \N__24914\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24908\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__24908\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__24905\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24899\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__24896\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24886\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24886\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24883\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24886\,
            I => \N__24880\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24883\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__24880\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24865\
        );

    \I__3463\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24865\
        );

    \I__3462\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24862\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24859\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24862\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__24859\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24848\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24848\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__24848\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__24833\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24821\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24821\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24821\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24815\,
            I => \N__24809\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24809\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24809\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__3442\ : CEMux
    port map (
            O => \N__24806\,
            I => \N__24785\
        );

    \I__3441\ : CEMux
    port map (
            O => \N__24805\,
            I => \N__24785\
        );

    \I__3440\ : CEMux
    port map (
            O => \N__24804\,
            I => \N__24785\
        );

    \I__3439\ : CEMux
    port map (
            O => \N__24803\,
            I => \N__24785\
        );

    \I__3438\ : CEMux
    port map (
            O => \N__24802\,
            I => \N__24785\
        );

    \I__3437\ : CEMux
    port map (
            O => \N__24801\,
            I => \N__24785\
        );

    \I__3436\ : CEMux
    port map (
            O => \N__24800\,
            I => \N__24785\
        );

    \I__3435\ : GlobalMux
    port map (
            O => \N__24785\,
            I => \N__24782\
        );

    \I__3434\ : gio2CtrlBuf
    port map (
            O => \N__24782\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__24779\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24770\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24775\,
            I => \N__24770\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__24770\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__24761\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df30\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__24758\,
            I => \N__24755\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24751\
        );

    \I__3424\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24748\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24751\,
            I => \N__24745\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24748\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__24745\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__24737\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__24734\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__3417\ : CascadeMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24725\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__3414\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24719\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__24719\,
            I => \N__24715\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24710\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__24715\,
            I => \N__24707\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24702\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24702\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__24710\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__24707\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24702\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__24689\,
            I => \N__24685\
        );

    \I__3402\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24682\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__24685\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__24682\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__24668\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__24665\,
            I => \N__24661\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__24664\,
            I => \N__24657\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24650\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24650\
        );

    \I__3391\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24650\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24650\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24644\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__24644\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__3386\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__24632\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24622\
        );

    \I__3382\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24622\
        );

    \I__3381\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24619\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__24622\,
            I => \N__24616\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__24619\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__24616\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3376\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24602\
        );

    \I__3375\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24602\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__24602\,
            I => \N__24598\
        );

    \I__3373\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24595\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__24598\,
            I => \N__24592\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__24595\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__24592\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__3369\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__24584\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__3367\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24575\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24575\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__24575\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__24572\,
            I => \N__24569\
        );

    \I__3363\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24563\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24563\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__24563\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__24560\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24554\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__24551\,
            I => \N__24548\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24545\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__3353\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__24536\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__24530\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__3349\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__24524\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__3347\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__24518\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__3345\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24506\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24506\
        );

    \I__3343\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24506\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__24506\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__24503\,
            I => \N__24498\
        );

    \I__3340\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24491\
        );

    \I__3339\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24491\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24491\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24487\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24484\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__24487\,
            I => \N__24481\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__24484\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__24481\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24467\
        );

    \I__3331\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24467\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24467\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24463\
        );

    \I__3328\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24460\
        );

    \I__3327\ : Span4Mux_v
    port map (
            O => \N__24463\,
            I => \N__24457\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__24460\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__24457\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24446\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__24443\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__24437\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24428\
        );

    \I__3317\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24428\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__24428\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24422\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__24422\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24410\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24410\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__24410\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__3309\ : InMux
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__24401\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24392\,
            I => \N__24389\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__24389\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__3301\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24380\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24371\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24371\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24367\
        );

    \I__3296\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24364\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__24367\,
            I => \N__24361\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__24364\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__24361\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24347\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24347\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24344\
        );

    \I__3288\ : Span4Mux_v
    port map (
            O => \N__24344\,
            I => \N__24340\
        );

    \I__3287\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24337\
        );

    \I__3286\ : Span4Mux_h
    port map (
            O => \N__24340\,
            I => \N__24334\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24337\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__24334\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__3283\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24326\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__24326\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__3281\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24317\
        );

    \I__3280\ : InMux
    port map (
            O => \N__24322\,
            I => \N__24317\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__24317\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__3277\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24305\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24305\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24305\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__24302\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__3272\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24293\,
            I => \N__24290\
        );

    \I__3270\ : Span4Mux_v
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__24287\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24278\
        );

    \I__3267\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24278\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__24278\,
            I => \N__24274\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24271\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__24274\,
            I => \N__24268\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__24271\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__24268\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24254\
        );

    \I__3259\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24254\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24250\
        );

    \I__3257\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24247\
        );

    \I__3256\ : Span4Mux_v
    port map (
            O => \N__24250\,
            I => \N__24244\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__24247\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__3254\ : Odrv4
    port map (
            O => \N__24244\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__3251\ : Span4Mux_v
    port map (
            O => \N__24233\,
            I => \N__24230\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__24230\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24221\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24214\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24225\,
            I => \N__24214\
        );

    \I__3246\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24214\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24221\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__24214\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3242\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24201\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24198\
        );

    \I__3240\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24195\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__24201\,
            I => \N__24190\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__24198\,
            I => \N__24190\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__24195\,
            I => \N__24183\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__24190\,
            I => \N__24183\
        );

    \I__3235\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24178\
        );

    \I__3234\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24178\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__24183\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__24178\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3231\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24170\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__24170\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__3229\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24164\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24164\,
            I => \N__24161\
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__24161\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__3225\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__24152\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24146\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__24146\,
            I => \N__24143\
        );

    \I__3221\ : Odrv12
    port map (
            O => \N__24143\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__3220\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__24137\,
            I => \N__24134\
        );

    \I__3218\ : Odrv12
    port map (
            O => \N__24134\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__24131\,
            I => \N__24127\
        );

    \I__3216\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24122\
        );

    \I__3215\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24122\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__24122\,
            I => \N__24118\
        );

    \I__3213\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24115\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__24118\,
            I => \N__24112\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__24115\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__24112\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__3209\ : InMux
    port map (
            O => \N__24107\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__3208\ : InMux
    port map (
            O => \N__24104\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24078\
        );

    \I__3206\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24078\
        );

    \I__3205\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24078\
        );

    \I__3204\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24078\
        );

    \I__3203\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24071\
        );

    \I__3202\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24071\
        );

    \I__3201\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24071\
        );

    \I__3200\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24062\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24062\
        );

    \I__3198\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24062\
        );

    \I__3197\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24062\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24090\,
            I => \N__24053\
        );

    \I__3195\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24053\
        );

    \I__3194\ : InMux
    port map (
            O => \N__24088\,
            I => \N__24053\
        );

    \I__3193\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24053\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24034\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__24071\,
            I => \N__24027\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__24062\,
            I => \N__24027\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24027\
        );

    \I__3188\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24020\
        );

    \I__3187\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24020\
        );

    \I__3186\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24020\
        );

    \I__3185\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24011\
        );

    \I__3184\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24011\
        );

    \I__3183\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24011\
        );

    \I__3182\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24011\
        );

    \I__3181\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24002\
        );

    \I__3180\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24002\
        );

    \I__3179\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24002\
        );

    \I__3178\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24002\
        );

    \I__3177\ : InMux
    port map (
            O => \N__24041\,
            I => \N__23993\
        );

    \I__3176\ : InMux
    port map (
            O => \N__24040\,
            I => \N__23993\
        );

    \I__3175\ : InMux
    port map (
            O => \N__24039\,
            I => \N__23993\
        );

    \I__3174\ : InMux
    port map (
            O => \N__24038\,
            I => \N__23993\
        );

    \I__3173\ : IoInMux
    port map (
            O => \N__24037\,
            I => \N__23990\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__24034\,
            I => \N__23977\
        );

    \I__3171\ : Span4Mux_v
    port map (
            O => \N__24027\,
            I => \N__23977\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__23977\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__23977\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23977\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23993\,
            I => \N__23977\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__23990\,
            I => \N__23974\
        );

    \I__3165\ : Span4Mux_v
    port map (
            O => \N__23977\,
            I => \N__23971\
        );

    \I__3164\ : Span12Mux_s8_v
    port map (
            O => \N__23974\,
            I => \N__23968\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__23971\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__3162\ : Odrv12
    port map (
            O => \N__23968\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23963\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__23954\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__3155\ : Span4Mux_v
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__23942\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__23939\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__23936\,
            I => \current_shift_inst.PI_CTRL.N_72_cascade_\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23930\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__23930\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23924\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23921\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23918\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23915\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23912\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23909\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23906\,
            I => \bfn_7_15_0_\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23903\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23900\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__23897\,
            I => \N__23894\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23890\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23887\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23881\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23881\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23878\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__23881\,
            I => \N__23875\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23878\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__23875\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23870\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23863\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23860\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23860\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__23857\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23852\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23845\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23842\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__23842\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__23839\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23834\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23828\,
            I => \N__23824\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23821\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__23824\,
            I => \N__23818\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__23821\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__23818\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23813\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23806\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23803\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23806\,
            I => \N__23800\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23803\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__23800\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23795\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23788\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23785\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__23788\,
            I => \N__23782\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__23785\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__3100\ : Odrv12
    port map (
            O => \N__23782\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23777\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23774\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23771\,
            I => \bfn_7_14_0_\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23761\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23761\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23758\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23761\,
            I => \N__23755\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23758\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3091\ : Odrv12
    port map (
            O => \N__23755\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23750\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__3088\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23738\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23738\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23734\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23737\,
            I => \N__23731\
        );

    \I__3084\ : Span4Mux_v
    port map (
            O => \N__23734\,
            I => \N__23728\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23731\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__23728\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23723\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23716\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23713\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23710\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23713\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__23710\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23705\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23698\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23695\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__23698\,
            I => \N__23692\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__23695\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__23692\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23687\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23681\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__23681\,
            I => \N__23677\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23674\
        );

    \I__3065\ : Span4Mux_v
    port map (
            O => \N__23677\,
            I => \N__23671\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__23674\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__23671\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__3062\ : InMux
    port map (
            O => \N__23666\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23656\
        );

    \I__3059\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23653\
        );

    \I__3058\ : Span4Mux_v
    port map (
            O => \N__23656\,
            I => \N__23650\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__23653\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__23650\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__3055\ : InMux
    port map (
            O => \N__23645\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__3054\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23638\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23635\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23632\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23635\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3050\ : Odrv12
    port map (
            O => \N__23632\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3049\ : InMux
    port map (
            O => \N__23627\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23620\
        );

    \I__3047\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23617\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__23620\,
            I => \N__23614\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23617\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3044\ : Odrv12
    port map (
            O => \N__23614\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3043\ : InMux
    port map (
            O => \N__23609\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23599\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23596\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__23599\,
            I => \N__23593\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__23596\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__23593\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3036\ : InMux
    port map (
            O => \N__23588\,
            I => \bfn_7_13_0_\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__23582\,
            I => \N__23578\
        );

    \I__3033\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23575\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__23578\,
            I => \N__23572\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__23575\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__3030\ : Odrv4
    port map (
            O => \N__23572\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23567\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__3028\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__23558\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__23555\,
            I => \N__23552\
        );

    \I__3024\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__23546\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23543\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23540\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23529\
        );

    \I__3017\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23526\
        );

    \I__3016\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23523\
        );

    \I__3015\ : Span4Mux_v
    port map (
            O => \N__23529\,
            I => \N__23518\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__23526\,
            I => \N__23518\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__23523\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__23518\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23509\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23506\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__23509\,
            I => \N__23503\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__23506\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__23503\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__3006\ : InMux
    port map (
            O => \N__23498\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__23489\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__23483\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23477\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23477\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__2997\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__23468\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__23465\,
            I => \N__23462\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23459\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__23447\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23441\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__2986\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__2984\ : Odrv12
    port map (
            O => \N__23432\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23420\
        );

    \I__2980\ : Odrv12
    port map (
            O => \N__23420\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__23417\,
            I => \N__23414\
        );

    \I__2978\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__23411\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__23408\,
            I => \N__23405\
        );

    \I__2975\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__23402\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__23399\,
            I => \N__23396\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__23393\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__23384\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__23375\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23369\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__23369\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__23360\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__2959\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23351\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__23351\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__2955\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__23339\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23333\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__23333\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__2949\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__23324\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__23312\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__2943\ : InMux
    port map (
            O => \N__23309\,
            I => \N__23303\
        );

    \I__2942\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23303\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__23303\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23291\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23291\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__23291\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__2936\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23284\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__23284\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__23281\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2932\ : InMux
    port map (
            O => \N__23276\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23269\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23269\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__23266\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23261\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__23255\,
            I => \N__23252\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__23252\,
            I => \N__23248\
        );

    \I__2923\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23245\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__23248\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23245\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2920\ : InMux
    port map (
            O => \N__23240\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__23237\,
            I => \N__23234\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23230\
        );

    \I__2917\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23227\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__23230\,
            I => \N__23222\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__23227\,
            I => \N__23222\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__23222\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2913\ : InMux
    port map (
            O => \N__23219\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2912\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23212\
        );

    \I__2911\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23209\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__23212\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__23209\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23204\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2907\ : InMux
    port map (
            O => \N__23201\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__2904\ : Span4Mux_s2_h
    port map (
            O => \N__23192\,
            I => \N__23184\
        );

    \I__2903\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23179\
        );

    \I__2902\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23179\
        );

    \I__2901\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23176\
        );

    \I__2900\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23173\
        );

    \I__2899\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23170\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__23184\,
            I => \N__23155\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__23179\,
            I => \N__23155\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23155\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__23173\,
            I => \N__23155\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23155\
        );

    \I__2893\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23152\
        );

    \I__2892\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23147\
        );

    \I__2891\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23147\
        );

    \I__2890\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23144\
        );

    \I__2889\ : Sp12to4
    port map (
            O => \N__23155\,
            I => \N__23137\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__23152\,
            I => \N__23137\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23137\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23134\
        );

    \I__2885\ : Span12Mux_v
    port map (
            O => \N__23137\,
            I => \N__23131\
        );

    \I__2884\ : Span12Mux_s5_h
    port map (
            O => \N__23134\,
            I => \N__23128\
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__23131\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2882\ : Odrv12
    port map (
            O => \N__23128\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__2880\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__2878\ : Odrv12
    port map (
            O => \N__23114\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2877\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23105\
        );

    \I__2876\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23105\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__23105\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23102\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__2872\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23092\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \N__23089\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23086\
        );

    \I__2869\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23083\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__23086\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__23083\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2866\ : InMux
    port map (
            O => \N__23078\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__2864\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23068\
        );

    \I__2863\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23065\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__23068\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__23065\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2860\ : InMux
    port map (
            O => \N__23060\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__23057\,
            I => \N__23053\
        );

    \I__2858\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23050\
        );

    \I__2857\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23047\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__23050\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__23047\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2854\ : InMux
    port map (
            O => \N__23042\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2853\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23035\
        );

    \I__2852\ : InMux
    port map (
            O => \N__23038\,
            I => \N__23032\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__23035\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__23032\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2849\ : InMux
    port map (
            O => \N__23027\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2848\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23021\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__23021\,
            I => \N__23017\
        );

    \I__2846\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23014\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__23017\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__23014\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2843\ : InMux
    port map (
            O => \N__23009\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2842\ : InMux
    port map (
            O => \N__23006\,
            I => \N__23000\
        );

    \I__2841\ : InMux
    port map (
            O => \N__23005\,
            I => \N__23000\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__23000\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22997\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22990\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22985\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22985\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22982\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__22982\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22979\,
            I => \bfn_5_18_0_\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22972\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22969\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22972\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__22969\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22964\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22958\,
            I => \N__22953\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22950\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22947\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__22953\,
            I => \N__22940\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22940\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22940\
        );

    \I__2820\ : Span4Mux_h
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__22937\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22934\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__22925\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22916\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22916\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22916\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2811\ : InMux
    port map (
            O => \N__22913\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22904\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22904\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__22904\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22901\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22895\,
            I => \N__22892\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__22892\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22886\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22886\,
            I => \N__22882\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__22882\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__22879\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22874\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__22865\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22856\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22856\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__22856\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2791\ : InMux
    port map (
            O => \N__22853\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22846\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22843\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22846\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22843\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22838\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2785\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22831\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22828\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22831\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__22828\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22823\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__22820\,
            I => \N__22817\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22813\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22810\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__22813\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22810\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22805\,
            I => \bfn_5_17_0_\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22799\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__22793\,
            I => \N__22790\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__22790\,
            I => \N__22787\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22787\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22784\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__22778\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__2763\ : Span4Mux_h
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__22766\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22763\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22754\,
            I => \N__22749\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22746\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22743\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__22749\,
            I => \N__22738\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22738\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__22743\,
            I => \N__22735\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__22738\,
            I => \N__22732\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__22735\,
            I => \N__22729\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__22732\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__22729\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22724\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22715\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__22712\,
            I => \N__22708\
        );

    \I__2743\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22704\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22698\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22698\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22695\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22692\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22698\,
            I => \N__22689\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__22695\,
            I => \N__22686\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__22692\,
            I => \N__22683\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__22689\,
            I => \N__22680\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__22686\,
            I => \N__22675\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__22683\,
            I => \N__22675\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__22680\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__22675\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22670\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2729\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__22661\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22651\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22648\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__22651\,
            I => \N__22642\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__22648\,
            I => \N__22642\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22639\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__22642\,
            I => \N__22636\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22633\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__22636\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__22633\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22628\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2715\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22622\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__22622\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22609\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22606\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__22609\,
            I => \N__22602\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22606\,
            I => \N__22599\
        );

    \I__2707\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22596\
        );

    \I__2706\ : Span4Mux_v
    port map (
            O => \N__22602\,
            I => \N__22593\
        );

    \I__2705\ : Span4Mux_h
    port map (
            O => \N__22599\,
            I => \N__22590\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__22596\,
            I => \N__22587\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__22593\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__22590\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__22587\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2700\ : InMux
    port map (
            O => \N__22580\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__22574\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22560\
        );

    \I__2694\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22557\
        );

    \I__2693\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22554\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__22560\,
            I => \N__22547\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__22557\,
            I => \N__22547\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22554\,
            I => \N__22547\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__22544\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22541\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22534\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22531\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22527\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22524\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22521\
        );

    \I__2681\ : Span4Mux_h
    port map (
            O => \N__22527\,
            I => \N__22518\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__22524\,
            I => \N__22513\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22513\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__22518\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__22513\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2676\ : InMux
    port map (
            O => \N__22508\,
            I => \bfn_5_16_0_\
        );

    \I__2675\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__22496\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2671\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__22490\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__2667\ : Odrv12
    port map (
            O => \N__22481\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__22478\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22471\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22468\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__22471\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__22468\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__2661\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22457\
        );

    \I__2660\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22457\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__22457\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__2658\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__22451\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__22448\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\
        );

    \I__2655\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__22439\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__22436\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__22433\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__2650\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__2648\ : Odrv12
    port map (
            O => \N__22424\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__2646\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__22415\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__22412\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22401\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__22408\,
            I => \N__22398\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22395\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22388\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22388\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22388\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__22401\,
            I => \N__22385\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22382\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22377\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22377\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__22385\,
            I => \N__22373\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22368\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__22377\,
            I => \N__22368\
        );

    \I__2630\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22365\
        );

    \I__2629\ : Span4Mux_v
    port map (
            O => \N__22373\,
            I => \N__22362\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__22368\,
            I => \N__22359\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22356\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__22362\,
            I => \current_shift_inst.PI_CTRL.N_164\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__22359\,
            I => \current_shift_inst.PI_CTRL.N_164\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__22356\,
            I => \current_shift_inst.PI_CTRL.N_164\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22346\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2620\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__22334\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__22322\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__22319\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__22313\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22307\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__22304\,
            I => \N__22300\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__22303\,
            I => \N__22297\
        );

    \I__2606\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22288\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22288\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22285\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22282\
        );

    \I__2602\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22276\
        );

    \I__2601\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22273\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__22288\,
            I => \N__22266\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__22285\,
            I => \N__22266\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__22282\,
            I => \N__22266\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22261\
        );

    \I__2596\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22261\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22258\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22253\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22253\
        );

    \I__2592\ : Span4Mux_s3_h
    port map (
            O => \N__22266\,
            I => \N__22250\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22247\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__22258\,
            I => \N__22244\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__22253\,
            I => \N__22241\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__22250\,
            I => \N__22236\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__22247\,
            I => \N__22236\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__22244\,
            I => \N__22233\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__22241\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__22236\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__22233\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2582\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__22223\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__22220\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__22214\,
            I => \current_shift_inst.PI_CTRL.N_71\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__22211\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__2576\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__22205\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__22199\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__2572\ : IoInMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2570\ : Span4Mux_s1_v
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2569\ : Sp12to4
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2568\ : Span12Mux_s10_h
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2567\ : Span12Mux_h
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2566\ : Span12Mux_v
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2565\ : Odrv12
    port map (
            O => \N__22175\,
            I => pwm_output_c
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__22166\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__2560\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__22157\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__22154\,
            I => \N__22151\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__22148\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__22139\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22133\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__2549\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22124\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__22121\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__22118\,
            I => \N__22111\
        );

    \I__2545\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22100\
        );

    \I__2544\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22100\
        );

    \I__2543\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22100\
        );

    \I__2542\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22100\
        );

    \I__2541\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22094\
        );

    \I__2540\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22089\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22089\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22086\
        );

    \I__2537\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22079\
        );

    \I__2536\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22079\
        );

    \I__2535\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22079\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__22094\,
            I => \N__22074\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22074\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__22086\,
            I => \N__22069\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__22079\,
            I => \N__22069\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__22074\,
            I => \N__22066\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__22069\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__22066\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__22061\,
            I => \N__22054\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__22060\,
            I => \N__22050\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__22059\,
            I => \N__22045\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__22058\,
            I => \N__22041\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__22057\,
            I => \N__22037\
        );

    \I__2522\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22032\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22032\
        );

    \I__2520\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22029\
        );

    \I__2519\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22020\
        );

    \I__2518\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22020\
        );

    \I__2517\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22020\
        );

    \I__2516\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22020\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22013\
        );

    \I__2514\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22013\
        );

    \I__2513\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22013\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__22032\,
            I => \N__21999\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__22029\,
            I => \N__21999\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__22020\,
            I => \N__21999\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__21999\
        );

    \I__2508\ : InMux
    port map (
            O => \N__22012\,
            I => \N__21979\
        );

    \I__2507\ : InMux
    port map (
            O => \N__22011\,
            I => \N__21979\
        );

    \I__2506\ : InMux
    port map (
            O => \N__22010\,
            I => \N__21972\
        );

    \I__2505\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21972\
        );

    \I__2504\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21972\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__21999\,
            I => \N__21969\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21951\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21951\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21951\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21951\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21951\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21951\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21951\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21951\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21936\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21936\
        );

    \I__2492\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21936\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21936\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21936\
        );

    \I__2489\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21936\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21936\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21931\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21931\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__21969\,
            I => \N__21928\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__21968\,
            I => \N__21925\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21917\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21936\,
            I => \N__21917\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__21931\,
            I => \N__21917\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__21928\,
            I => \N__21914\
        );

    \I__2479\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21911\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21908\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__21917\,
            I => \N__21905\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__21914\,
            I => \N_19_1\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__21911\,
            I => \N_19_1\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N_19_1\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__21905\,
            I => \N_19_1\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21890\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1\
        );

    \I__2469\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21872\
        );

    \I__2468\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21872\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21872\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21872\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21865\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21865\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21865\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21857\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21857\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21850\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21863\,
            I => \N__21850\
        );

    \I__2458\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21850\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__21857\,
            I => \N__21845\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21845\
        );

    \I__2455\ : Span4Mux_v
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__21842\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__21830\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__21827\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__21815\,
            I => \N__21811\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21808\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__21811\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21808\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__21800\,
            I => \N__21796\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21792\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__21796\,
            I => \N__21789\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21786\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__21792\,
            I => \N__21781\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__21789\,
            I => \N__21781\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21786\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__21781\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21773\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__21764\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21754\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21750\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__21754\,
            I => \N__21747\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21744\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21750\,
            I => \N__21741\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__21747\,
            I => \N__21738\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21744\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2419\ : Odrv12
    port map (
            O => \N__21741\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__21738\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__21728\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__2414\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21719\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__2412\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21712\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21709\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21706\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__21709\,
            I => \N__21703\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__21706\,
            I => \N__21699\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__21703\,
            I => \N__21696\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21693\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__21699\,
            I => \N__21690\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__21696\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__21693\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__21690\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2401\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21680\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__21668\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__2395\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21661\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21658\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21655\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21658\,
            I => \N__21651\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__21655\,
            I => \N__21648\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21645\
        );

    \I__2389\ : Span12Mux_h
    port map (
            O => \N__21651\,
            I => \N__21642\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__21648\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__21645\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__21642\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__21632\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21625\
        );

    \I__2382\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21622\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__21625\,
            I => \N__21619\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__21622\,
            I => \N__21615\
        );

    \I__2379\ : Span4Mux_h
    port map (
            O => \N__21619\,
            I => \N__21612\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21609\
        );

    \I__2377\ : Span4Mux_h
    port map (
            O => \N__21615\,
            I => \N__21606\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__21612\,
            I => \N__21603\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21609\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__21606\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__21603\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2372\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21593\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__21593\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2370\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__21587\,
            I => \N__21583\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21579\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__21583\,
            I => \N__21576\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21573\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__21579\,
            I => \N__21566\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__21576\,
            I => \N__21566\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21566\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__21566\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21560\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21554\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21554\,
            I => \N__21551\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__21551\,
            I => \N__21546\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21543\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21540\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__21546\,
            I => \N__21535\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__21543\,
            I => \N__21535\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21540\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__21535\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__21527\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2348\ : InMux
    port map (
            O => \N__21524\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2347\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21503\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21503\
        );

    \I__2345\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21503\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21503\
        );

    \I__2343\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21494\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21494\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21494\
        );

    \I__2340\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21494\
        );

    \I__2339\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21489\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21489\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21503\,
            I => \N__21484\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21484\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__21489\,
            I => \N__21481\
        );

    \I__2334\ : Span4Mux_s3_h
    port map (
            O => \N__21484\,
            I => \N__21478\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__21481\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__21478\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21473\,
            I => \N__21467\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21460\
        );

    \I__2329\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21460\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21460\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21457\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__21460\,
            I => \N__21454\
        );

    \I__2325\ : Span4Mux_s3_h
    port map (
            O => \N__21457\,
            I => \N__21450\
        );

    \I__2324\ : Span4Mux_s3_h
    port map (
            O => \N__21454\,
            I => \N__21447\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21444\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__21450\,
            I => \current_shift_inst.PI_CTRL.N_144\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__21447\,
            I => \current_shift_inst.PI_CTRL.N_144\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__21444\,
            I => \current_shift_inst.PI_CTRL.N_144\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__21431\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1\
        );

    \I__2316\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__21422\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__21419\,
            I => \N__21416\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__21413\,
            I => \current_shift_inst.PI_CTRL.N_146\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__2307\ : Span4Mux_h
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__21398\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__21389\,
            I => \N__21386\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__21386\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21376\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21372\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__21376\,
            I => \N__21369\
        );

    \I__2297\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21366\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21363\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__21369\,
            I => \N__21360\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__21366\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__21363\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__21360\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__21350\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__21338\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21328\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21324\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__21328\,
            I => \N__21321\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21318\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__21324\,
            I => \N__21315\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__21321\,
            I => \N__21312\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21318\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__21315\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__21312\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2275\ : InMux
    port map (
            O => \N__21305\,
            I => \N__21302\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21302\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__21299\,
            I => \N__21296\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__21293\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__2270\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21287\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21284\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__21284\,
            I => \N__21279\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21276\
        );

    \I__2266\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21273\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__21279\,
            I => \N__21268\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__21276\,
            I => \N__21268\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21273\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__21268\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2261\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__21260\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__21251\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__2256\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21245\,
            I => \N__21242\
        );

    \I__2254\ : Odrv12
    port map (
            O => \N__21242\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__21239\,
            I => \N__21235\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__21238\,
            I => \N__21231\
        );

    \I__2251\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21227\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21224\
        );

    \I__2249\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21221\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__21230\,
            I => \N__21215\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21227\,
            I => \N__21211\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21208\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21205\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__21220\,
            I => \N__21200\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__21219\,
            I => \N__21197\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21192\
        );

    \I__2241\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21189\
        );

    \I__2240\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21186\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__21211\,
            I => \N__21183\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__21208\,
            I => \N__21178\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__21205\,
            I => \N__21178\
        );

    \I__2236\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21165\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21165\
        );

    \I__2234\ : InMux
    port map (
            O => \N__21200\,
            I => \N__21165\
        );

    \I__2233\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21165\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21165\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21165\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21158\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__21189\,
            I => \N__21158\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21158\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__21183\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__21178\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__21165\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2224\ : Odrv12
    port map (
            O => \N__21158\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21149\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__2221\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21136\
        );

    \I__2219\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21133\
        );

    \I__2218\ : Sp12to4
    port map (
            O => \N__21136\,
            I => \N__21128\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21128\
        );

    \I__2216\ : Odrv12
    port map (
            O => \N__21128\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__2215\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21121\
        );

    \I__2214\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21117\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21114\
        );

    \I__2212\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21111\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__21117\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__21114\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__21111\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2208\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21097\
        );

    \I__2206\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21094\
        );

    \I__2205\ : Sp12to4
    port map (
            O => \N__21097\,
            I => \N__21089\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21089\
        );

    \I__2203\ : Odrv12
    port map (
            O => \N__21089\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__2201\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21078\
        );

    \I__2200\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21075\
        );

    \I__2199\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21072\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__21078\,
            I => \N__21069\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__21075\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__21072\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__21069\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2194\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21058\
        );

    \I__2193\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21055\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21052\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__21055\,
            I => \N__21049\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__21052\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__21049\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\
        );

    \I__2188\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__21041\,
            I => \N__21037\
        );

    \I__2186\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21033\
        );

    \I__2185\ : Span4Mux_s2_h
    port map (
            O => \N__21037\,
            I => \N__21030\
        );

    \I__2184\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21027\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__21033\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__21030\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__21027\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2180\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21014\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__21014\,
            I => un7_start_stop_0_a2
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__21011\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__21008\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__2175\ : InMux
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__21002\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__20999\,
            I => \N__20996\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__20990\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__20984\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20981\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20975\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__20969\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__20966\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__20960\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20957\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20951\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20948\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20942\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20936\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20933\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20927\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20924\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20918\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20915\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20909\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20906\,
            I => \bfn_2_18_0_\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__20897\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__20888\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__20879\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__20870\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20867\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__20861\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20855\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__20843\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20840\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__20831\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20828\,
            I => \bfn_2_15_0_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__20819\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__20810\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__20801\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\
        );

    \I__2106\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__20795\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__20789\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20783\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20783\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20777\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__20774\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20766\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20761\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20761\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20766\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20761\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20753\,
            I => \N__20749\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20746\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20740\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__20743\,
            I => \N__20737\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__20740\,
            I => \N__20734\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__20737\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__20734\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__20720\,
            I => \pwm_generator_inst.O_12\
        );

    \I__2079\ : InMux
    port map (
            O => \N__20717\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20708\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__20705\,
            I => \pwm_generator_inst.O_13\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__20696\,
            I => \N__20692\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20689\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__20692\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20689\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20684\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__2067\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__20672\,
            I => \pwm_generator_inst.O_14\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20662\
        );

    \I__2061\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20659\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__20662\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__20659\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2058\ : InMux
    port map (
            O => \N__20654\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20648\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__2055\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__20642\,
            I => \N__20638\
        );

    \I__2053\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20635\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__20638\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__20635\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2050\ : InMux
    port map (
            O => \N__20630\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__20621\,
            I => \N__20618\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__20618\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\
        );

    \I__2045\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20608\
        );

    \I__2043\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20605\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__20608\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__20605\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20600\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__20594\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20591\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__2036\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20580\
        );

    \I__2034\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20575\
        );

    \I__2033\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20575\
        );

    \I__2032\ : Span4Mux_s2_h
    port map (
            O => \N__20580\,
            I => \N__20572\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__20575\,
            I => pwm_duty_input_6
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__20572\,
            I => pwm_duty_input_6
        );

    \I__2029\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20560\
        );

    \I__2028\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20560\
        );

    \I__2027\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20557\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__20560\,
            I => pwm_duty_input_8
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__20557\,
            I => pwm_duty_input_8
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__20552\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20545\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__20548\,
            I => \N__20541\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__20545\,
            I => \N__20538\
        );

    \I__2020\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20533\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20533\
        );

    \I__2018\ : Span4Mux_s1_h
    port map (
            O => \N__20538\,
            I => \N__20530\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__20533\,
            I => pwm_duty_input_9
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__20530\,
            I => pwm_duty_input_9
        );

    \I__2015\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20522\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20517\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20514\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20511\
        );

    \I__2011\ : Span4Mux_s1_h
    port map (
            O => \N__20517\,
            I => \N__20508\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__20514\,
            I => pwm_duty_input_3
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__20511\,
            I => pwm_duty_input_3
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__20508\,
            I => pwm_duty_input_3
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__20501\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20490\
        );

    \I__2004\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20487\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20484\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__20490\,
            I => \N__20481\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__20487\,
            I => pwm_duty_input_4
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__20484\,
            I => pwm_duty_input_4
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__20481\,
            I => pwm_duty_input_4
        );

    \I__1998\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__20471\,
            I => \N__20467\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20464\
        );

    \I__1995\ : Span4Mux_s1_h
    port map (
            O => \N__20467\,
            I => \N__20461\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20464\,
            I => pwm_duty_input_0
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__20461\,
            I => pwm_duty_input_0
        );

    \I__1992\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20452\
        );

    \I__1991\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__20452\,
            I => pwm_duty_input_1
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__20449\,
            I => pwm_duty_input_1
        );

    \I__1988\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20440\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20437\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__20440\,
            I => pwm_duty_input_2
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20437\,
            I => pwm_duty_input_2
        );

    \I__1984\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__20429\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__1982\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__20420\,
            I => \current_shift_inst.PI_CTRL.N_140\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__20411\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__20408\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__20405\,
            I => \N__20400\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__20404\,
            I => \N__20397\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__20403\,
            I => \N__20394\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20400\,
            I => \N__20391\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20397\,
            I => \N__20386\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20386\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20391\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__20386\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1967\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20372\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20372\
        );

    \I__1965\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20372\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__20369\,
            I => \current_shift_inst.PI_CTRL.N_145\
        );

    \I__1962\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20358\
        );

    \I__1960\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20355\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20352\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__20358\,
            I => \N__20349\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20355\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__20352\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__20349\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__1953\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__1951\ : Odrv12
    port map (
            O => \N__20333\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__1950\ : InMux
    port map (
            O => \N__20330\,
            I => \bfn_1_21_0_\
        );

    \I__1949\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__1947\ : Odrv12
    port map (
            O => \N__20321\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__1946\ : InMux
    port map (
            O => \N__20318\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__20309\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__1942\ : InMux
    port map (
            O => \N__20306\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__1941\ : InMux
    port map (
            O => \N__20303\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__1940\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N_42_i_i\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__20291\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20281\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20281\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20278\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20281\,
            I => pwm_duty_input_7
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20278\,
            I => pwm_duty_input_7
        );

    \I__1931\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20269\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__20272\,
            I => \N__20266\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20262\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20259\
        );

    \I__1927\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20256\
        );

    \I__1926\ : Span4Mux_s1_h
    port map (
            O => \N__20262\,
            I => \N__20253\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20259\,
            I => pwm_duty_input_5
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20256\,
            I => pwm_duty_input_5
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__20253\,
            I => pwm_duty_input_5
        );

    \I__1922\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__1920\ : Span4Mux_v
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__20234\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1917\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__20228\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__1913\ : Span12Mux_h
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__20216\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1911\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__20210\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__1909\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20204\,
            I => \N__20200\
        );

    \I__1907\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__20200\,
            I => \N__20194\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20197\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__20194\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__20183\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__1900\ : InMux
    port map (
            O => \N__20180\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__1899\ : InMux
    port map (
            O => \N__20177\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__1898\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__20171\,
            I => \N__20168\
        );

    \I__1896\ : Odrv12
    port map (
            O => \N__20168\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__1895\ : InMux
    port map (
            O => \N__20165\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20157\
        );

    \I__1893\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20154\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20151\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__20157\,
            I => \N__20148\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__20154\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__20151\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__1888\ : Odrv12
    port map (
            O => \N__20148\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__20138\,
            I => \N__20135\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__20135\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__1884\ : InMux
    port map (
            O => \N__20132\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__1883\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20124\
        );

    \I__1882\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20121\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20118\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__20124\,
            I => \N__20115\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__20121\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__20118\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__1877\ : Odrv12
    port map (
            O => \N__20115\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__1876\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__20096\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__1871\ : InMux
    port map (
            O => \N__20093\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \N__20086\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__20089\,
            I => \N__20082\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20079\
        );

    \I__1867\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20076\
        );

    \I__1866\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20073\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__20079\,
            I => \N__20070\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__20076\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__20073\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__20070\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__1861\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__1859\ : Odrv12
    port map (
            O => \N__20057\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__1858\ : InMux
    port map (
            O => \N__20054\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__1857\ : InMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__20039\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1852\ : InMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__20033\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__1850\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__1848\ : Span12Mux_h
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__1847\ : Odrv12
    port map (
            O => \N__20021\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1846\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__20015\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__1844\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__20009\,
            I => \N__20006\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__20000\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__19994\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__19976\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__19970\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__1829\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__19955\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__19949\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__1820\ : Span4Mux_v
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__19934\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1817\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19928\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__19913\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19907\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__19892\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__19886\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19877\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19877\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__19871\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__19868\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10_cascade_\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__19850\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19847\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__1787\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__1783\ : Odrv4
    port map (
            O => \N__19829\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19826\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19808\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19805\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__1774\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19796\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19796\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19793\,
            I => \N__19784\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19777\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19777\
        );

    \I__1768\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19777\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19770\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19770\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19770\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__19784\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__19777\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__19770\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__19754\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19751\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__1754\ : Span12Mux_v
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__1753\ : Odrv12
    port map (
            O => \N__19739\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__1752\ : InMux
    port map (
            O => \N__19736\,
            I => \bfn_1_15_0_\
        );

    \I__1751\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__19721\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__19712\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19709\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__19694\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19685\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__1734\ : InMux
    port map (
            O => \N__19682\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__1733\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__19667\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__1727\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__19658\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__1725\ : InMux
    port map (
            O => \N__19655\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__19640\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19631\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__1716\ : InMux
    port map (
            O => \N__19628\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__1715\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__1713\ : Span12Mux_h
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__19616\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1710\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__19601\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__1706\ : InMux
    port map (
            O => \N__19598\,
            I => \bfn_1_14_0_\
        );

    \I__1705\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__19592\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1702\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__19574\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19571\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__19553\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__1690\ : InMux
    port map (
            O => \N__19550\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__19532\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__1683\ : InMux
    port map (
            O => \N__19529\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__1680\ : Span12Mux_h
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__19517\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__1677\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__19502\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__19487\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19478\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19475\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__1662\ : Span4Mux_v
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__19460\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__19451\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__1656\ : InMux
    port map (
            O => \N__19448\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__19436\,
            I => \N__19433\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__19433\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__1649\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__19424\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__1647\ : InMux
    port map (
            O => \N__19421\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19418\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__1645\ : InMux
    port map (
            O => \N__19415\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__1644\ : InMux
    port map (
            O => \N__19412\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19409\,
            I => \bfn_1_10_0_\
        );

    \I__1642\ : InMux
    port map (
            O => \N__19406\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__1641\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__19400\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__1639\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19391\
        );

    \I__1638\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19391\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__19391\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1636\ : InMux
    port map (
            O => \N__19388\,
            I => \bfn_1_9_0_\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19385\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__1634\ : InMux
    port map (
            O => \N__19382\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__1633\ : InMux
    port map (
            O => \N__19379\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__1632\ : InMux
    port map (
            O => \N__19376\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__1631\ : IoInMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__1629\ : Span4Mux_s3_v
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1628\ : Span4Mux_h
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__1627\ : Sp12to4
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__1626\ : Span12Mux_s9_v
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1625\ : Span12Mux_v
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1624\ : Odrv12
    port map (
            O => \N__19352\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1623\ : IoInMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__1621\ : IoSpan4Mux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__1620\ : IoSpan4Mux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__19337\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_18_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_7_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_12_14_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19373\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19349\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35582\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_167_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24037\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__37436\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__45040\,
            CLKHFEN => \N__45044\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__45088\,
            RGB2PWM => \N__20300\,
            RGB1 => rgb_g_wire,
            CURREN => \N__45045\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__21020\,
            RGB0PWM => \N__48683\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23198\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49148\,
            ce => 'H',
            sr => \N__48597\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__19397\,
            in1 => \N__19403\,
            in2 => \N__21968\,
            in3 => \N__19801\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__19396\,
            in1 => \N__21924\,
            in2 => \_gnd_net_\,
            in3 => \N__19802\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21518\,
            in1 => \N__21375\,
            in2 => \_gnd_net_\,
            in3 => \N__19388\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21514\,
            in1 => \N__21327\,
            in2 => \_gnd_net_\,
            in3 => \N__19385\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_2_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21519\,
            in1 => \N__21282\,
            in2 => \_gnd_net_\,
            in3 => \N__19382\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_3_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21515\,
            in1 => \N__21795\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_4_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__21753\,
            in2 => \_gnd_net_\,
            in3 => \N__19376\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_5_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21516\,
            in1 => \N__21702\,
            in2 => \_gnd_net_\,
            in3 => \N__19418\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_6_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21521\,
            in1 => \N__21654\,
            in2 => \_gnd_net_\,
            in3 => \N__19415\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_7_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21517\,
            in1 => \N__21618\,
            in2 => \_gnd_net_\,
            in3 => \N__19412\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__49147\,
            ce => 'H',
            sr => \N__48629\
        );

    \pwm_generator_inst.counter_8_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21513\,
            in1 => \N__21586\,
            in2 => \_gnd_net_\,
            in3 => \N__19409\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__49146\,
            ce => 'H',
            sr => \N__48636\
        );

    \pwm_generator_inst.counter_9_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21549\,
            in1 => \N__21512\,
            in2 => \_gnd_net_\,
            in3 => \N__19406\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => 'H',
            sr => \N__48636\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__22404\,
            in1 => \N__22711\,
            in2 => \N__21824\,
            in3 => \N__20426\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => 'H',
            sr => \N__48636\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111010"
        )
    port map (
            in0 => \N__22658\,
            in1 => \N__22405\,
            in2 => \N__22303\,
            in3 => \N__23190\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => 'H',
            sr => \N__48636\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111010"
        )
    port map (
            in0 => \N__22961\,
            in1 => \N__22406\,
            in2 => \N__22304\,
            in3 => \N__23191\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => 'H',
            sr => \N__48636\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__22295\,
            in1 => \N__20417\,
            in2 => \N__22760\,
            in3 => \N__21473\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => 'H',
            sr => \N__48636\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__21471\,
            in1 => \N__22775\,
            in2 => \N__20404\,
            in3 => \N__20381\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49144\,
            ce => 'H',
            sr => \N__48639\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20379\,
            in1 => \N__22505\,
            in2 => \N__20405\,
            in3 => \N__21472\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49144\,
            ce => 'H',
            sr => \N__48639\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__23189\,
            in1 => \N__22294\,
            in2 => \N__22571\,
            in3 => \N__22407\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49144\,
            ce => 'H',
            sr => \N__48639\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__21470\,
            in1 => \N__22796\,
            in2 => \N__20403\,
            in3 => \N__20380\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49144\,
            ce => 'H',
            sr => \N__48639\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__22537\,
            in1 => \N__22293\,
            in2 => \N__22408\,
            in3 => \N__23187\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49141\,
            ce => 'H',
            sr => \N__48643\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19526\,
            in2 => \N__19514\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19499\,
            in2 => \N__19484\,
            in3 => \N__19475\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19472\,
            in2 => \N__19457\,
            in3 => \N__19448\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19445\,
            in2 => \N__19430\,
            in3 => \N__19421\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19733\,
            in2 => \N__19718\,
            in3 => \N__19709\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19706\,
            in2 => \N__19691\,
            in3 => \N__19682\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19679\,
            in2 => \N__19664\,
            in3 => \N__19655\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19652\,
            in2 => \N__19637\,
            in3 => \N__19628\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19625\,
            in2 => \N__19613\,
            in3 => \N__19598\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19595\,
            in2 => \N__19589\,
            in3 => \N__19571\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19787\,
            in2 => \N__19568\,
            in3 => \N__19550\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19790\,
            in2 => \N__19547\,
            in3 => \N__19529\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19788\,
            in2 => \N__19865\,
            in3 => \N__19847\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19791\,
            in2 => \N__19844\,
            in3 => \N__19826\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19789\,
            in2 => \N__19823\,
            in3 => \N__19805\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19792\,
            in2 => \N__19763\,
            in3 => \N__19751\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19748\,
            in1 => \N__20864\,
            in2 => \_gnd_net_\,
            in3 => \N__19736\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20085\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20641\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27628\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20665\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20695\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20362\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20611\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19882\,
            in2 => \_gnd_net_\,
            in3 => \N__20203\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__19883\,
            in1 => \N__21195\,
            in2 => \N__19868\,
            in3 => \N__20189\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20702\,
            in1 => \N__20141\,
            in2 => \N__21219\,
            in3 => \N__20160\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__21125\,
            in1 => \N__21196\,
            in2 => \N__21146\,
            in3 => \N__20174\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20669\,
            in1 => \N__20108\,
            in2 => \N__21220\,
            in3 => \N__20127\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__20615\,
            in1 => \N__21204\,
            in2 => \N__20342\,
            in3 => \N__20361\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__21203\,
            in1 => \N__20645\,
            in2 => \N__20089\,
            in3 => \N__20063\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21062\,
            in1 => \N__20327\,
            in2 => \N__21230\,
            in3 => \N__21044\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__21104\,
            in1 => \N__21218\,
            in2 => \N__21086\,
            in3 => \N__20315\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20036\,
            in2 => \_gnd_net_\,
            in3 => \N__20051\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20018\,
            in2 => \_gnd_net_\,
            in3 => \N__20030\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19997\,
            in2 => \_gnd_net_\,
            in3 => \N__20012\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19973\,
            in2 => \_gnd_net_\,
            in3 => \N__19991\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19952\,
            in2 => \_gnd_net_\,
            in3 => \N__19967\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19931\,
            in2 => \_gnd_net_\,
            in3 => \N__19946\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19910\,
            in2 => \_gnd_net_\,
            in3 => \N__19925\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19889\,
            in2 => \_gnd_net_\,
            in3 => \N__19904\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20231\,
            in2 => \_gnd_net_\,
            in3 => \N__20246\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20213\,
            in2 => \_gnd_net_\,
            in3 => \N__20225\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20207\,
            in2 => \_gnd_net_\,
            in3 => \N__20180\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__21214\,
            in1 => \N__20756\,
            in2 => \_gnd_net_\,
            in3 => \N__20177\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21120\,
            in2 => \_gnd_net_\,
            in3 => \N__20165\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20162\,
            in2 => \_gnd_net_\,
            in3 => \N__20132\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20129\,
            in2 => \_gnd_net_\,
            in3 => \N__20093\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20090\,
            in3 => \N__20054\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20366\,
            in2 => \_gnd_net_\,
            in3 => \N__20330\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21036\,
            in2 => \_gnd_net_\,
            in3 => \N__20318\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21081\,
            in2 => \_gnd_net_\,
            in3 => \N__20306\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20303\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.N_42_i_i_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35066\,
            in2 => \_gnd_net_\,
            in3 => \N__48682\,
            lcout => \N_42_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20521\,
            in1 => \N__20494\,
            in2 => \N__20272\,
            in3 => \N__20294\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__23188\,
            in1 => \N__22296\,
            in2 => \N__22619\,
            in3 => \N__22409\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => 'H',
            sr => \N__48630\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20566\,
            in1 => \N__20583\,
            in2 => \N__20548\,
            in3 => \N__20288\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20287\,
            in2 => \_gnd_net_\,
            in3 => \N__20265\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20584\,
            in1 => \N__20567\,
            in2 => \N__20552\,
            in3 => \N__20544\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__20432\,
            in1 => \N__20520\,
            in2 => \N__20501\,
            in3 => \N__20493\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20470\,
            in1 => \N__20456\,
            in2 => \_gnd_net_\,
            in3 => \N__20444\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__20770\,
            in1 => \N__23168\,
            in2 => \N__22712\,
            in3 => \N__22280\,
            lcout => \current_shift_inst.PI_CTRL.N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__23167\,
            in1 => \N__22707\,
            in2 => \_gnd_net_\,
            in3 => \N__20769\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__22753\,
            in1 => \N__22281\,
            in2 => \N__20408\,
            in3 => \N__21453\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__23169\,
            in1 => \N__20771\,
            in2 => \_gnd_net_\,
            in3 => \N__22279\,
            lcout => \current_shift_inst.PI_CTRL.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22956\,
            in2 => \_gnd_net_\,
            in3 => \N__22654\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22564\,
            in1 => \N__22612\,
            in2 => \N__20774\,
            in3 => \N__22538\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20752\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20729\,
            in2 => \_gnd_net_\,
            in3 => \N__20717\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20714\,
            in2 => \_gnd_net_\,
            in3 => \N__20684\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20681\,
            in2 => \_gnd_net_\,
            in3 => \N__20654\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20651\,
            in2 => \_gnd_net_\,
            in3 => \N__20630\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44868\,
            in2 => \N__20627\,
            in3 => \N__20600\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20597\,
            in2 => \N__44924\,
            in3 => \N__20591\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44872\,
            in2 => \N__20852\,
            in3 => \N__20840\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20837\,
            in2 => \_gnd_net_\,
            in3 => \N__20828\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20825\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20816\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20807\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20798\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20792\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20786\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20780\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20903\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20894\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20885\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20876\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20867\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__22109\,
            in1 => \N__20987\,
            in2 => \N__22057\,
            in3 => \N__21881\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__21882\,
            in1 => \N__22040\,
            in2 => \N__22118\,
            in3 => \N__20972\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__22110\,
            in1 => \N__20939\,
            in2 => \N__22058\,
            in3 => \N__21883\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20858\,
            in2 => \N__21238\,
            in3 => \N__21234\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31\,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20999\,
            in3 => \N__20981\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20978\,
            in2 => \_gnd_net_\,
            in3 => \N__20966\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20963\,
            in2 => \_gnd_net_\,
            in3 => \N__20957\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20954\,
            in2 => \_gnd_net_\,
            in3 => \N__20948\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20945\,
            in2 => \_gnd_net_\,
            in3 => \N__20933\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20930\,
            in2 => \_gnd_net_\,
            in3 => \N__20924\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20921\,
            in2 => \_gnd_net_\,
            in3 => \N__20915\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20912\,
            in2 => \_gnd_net_\,
            in3 => \N__20906\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__21257\,
            in1 => \N__21248\,
            in2 => \N__21239\,
            in3 => \N__21149\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21139\,
            in2 => \_gnd_net_\,
            in3 => \N__21124\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21082\,
            in2 => \_gnd_net_\,
            in3 => \N__21100\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21061\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un7_start_stop_0_a2_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35065\,
            in2 => \_gnd_net_\,
            in3 => \N__48681\,
            lcout => un7_start_stop_0_a2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21283\,
            in2 => \_gnd_net_\,
            in3 => \N__21379\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__21757\,
            in1 => \N__21799\,
            in2 => \N__21011\,
            in3 => \N__21331\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21550\,
            in1 => \N__21582\,
            in2 => \_gnd_net_\,
            in3 => \N__21628\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21665\,
            in1 => \N__21715\,
            in2 => \N__21008\,
            in3 => \N__21005\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__23166\,
            in1 => \N__21814\,
            in2 => \N__21419\,
            in3 => \N__22376\,
            lcout => \current_shift_inst.PI_CTRL.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21863\,
            in1 => \N__22099\,
            in2 => \N__22061\,
            in3 => \N__21437\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__22097\,
            in1 => \N__21428\,
            in2 => \N__22060\,
            in3 => \N__21862\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22703\,
            in2 => \_gnd_net_\,
            in3 => \N__22752\,
            lcout => \current_shift_inst.PI_CTRL.N_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__22098\,
            in1 => \N__22053\,
            in2 => \N__21410\,
            in3 => \N__21864\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21353\,
            in2 => \N__21395\,
            in3 => \N__21383\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21305\,
            in2 => \N__21347\,
            in3 => \N__21335\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21263\,
            in2 => \N__21299\,
            in3 => \N__21290\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21776\,
            in2 => \N__21839\,
            in3 => \N__21803\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21731\,
            in2 => \N__21770\,
            in3 => \N__21761\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21683\,
            in2 => \N__21725\,
            in3 => \N__21716\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21635\,
            in2 => \N__21677\,
            in3 => \N__21664\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21596\,
            in2 => \N__22130\,
            in3 => \N__21629\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21563\,
            in2 => \N__22145\,
            in3 => \N__21590\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21530\,
            in2 => \N__22163\,
            in3 => \N__21557\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21524\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49109\,
            ce => 'H',
            sr => \N__48652\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__22117\,
            in1 => \N__21887\,
            in2 => \N__22172\,
            in3 => \N__22049\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__22116\,
            in1 => \N__22048\,
            in2 => \N__22154\,
            in3 => \N__21886\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__21885\,
            in1 => \N__22115\,
            in2 => \N__22059\,
            in3 => \N__22136\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27422\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__22114\,
            in1 => \N__22044\,
            in2 => \N__21896\,
            in3 => \N__21884\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__22530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22647\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22605\,
            in1 => \N__22563\,
            in2 => \N__21827\,
            in3 => \N__22957\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22487\,
            in1 => \N__22430\,
            in2 => \N__22343\,
            in3 => \N__22328\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28301\,
            in1 => \N__30095\,
            in2 => \N__27430\,
            in3 => \N__32032\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001011"
        )
    port map (
            in0 => \N__22202\,
            in1 => \N__25018\,
            in2 => \N__27206\,
            in3 => \N__22208\,
            lcout => \current_shift_inst.PI_CTRL.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29766\,
            in1 => \N__27813\,
            in2 => \N__29834\,
            in3 => \N__29914\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22226\,
            in1 => \N__22445\,
            in2 => \N__22220\,
            in3 => \N__22217\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24205\,
            in2 => \_gnd_net_\,
            in3 => \N__27153\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__27862\,
            in1 => \N__31856\,
            in2 => \N__22211\,
            in3 => \N__27529\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__27259\,
            in1 => \N__27104\,
            in2 => \_gnd_net_\,
            in3 => \N__26959\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22885\,
            in2 => \_gnd_net_\,
            in3 => \N__22921\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22993\,
            in1 => \N__23006\,
            in2 => \N__23237\,
            in3 => \N__23038\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23258\,
            in1 => \N__22909\,
            in2 => \N__22421\,
            in3 => \N__22418\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22310\,
            in1 => \N__22349\,
            in2 => \N__22412\,
            in3 => \N__22316\,
            lcout => \current_shift_inst.PI_CTRL.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23071\,
            in1 => \N__22849\,
            in2 => \N__23057\,
            in3 => \N__22861\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22862\,
            in1 => \N__22850\,
            in2 => \N__22994\,
            in3 => \N__23005\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23233\,
            in1 => \N__22922\,
            in2 => \N__22820\,
            in3 => \N__22835\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22910\,
            in1 => \N__22889\,
            in2 => \N__22331\,
            in3 => \N__22454\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22816\,
            in2 => \_gnd_net_\,
            in3 => \N__22834\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23024\,
            in1 => \N__22975\,
            in2 => \N__22319\,
            in3 => \N__23287\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23272\,
            in1 => \N__23111\,
            in2 => \N__23099\,
            in3 => \N__23216\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__23110\,
            in1 => \_gnd_net_\,
            in2 => \N__23095\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27692\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27371\,
            in1 => \N__27693\,
            in2 => \N__41284\,
            in3 => \N__27744\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24140\,
            in1 => \N__24149\,
            in2 => \N__22448\,
            in3 => \N__24167\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28293\,
            in2 => \_gnd_net_\,
            in3 => \N__27423\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22493\,
            in1 => \N__25498\,
            in2 => \N__22436\,
            in3 => \N__30089\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23215\,
            in2 => \_gnd_net_\,
            in3 => \N__23273\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23251\,
            in1 => \N__23020\,
            in2 => \N__22433\,
            in3 => \N__23039\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27365\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29910\,
            in1 => \N__29756\,
            in2 => \N__29835\,
            in3 => \N__27809\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23056\,
            in1 => \N__22976\,
            in2 => \N__23075\,
            in3 => \N__23288\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26795\,
            in2 => \_gnd_net_\,
            in3 => \N__24722\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__26743\,
            in1 => \N__24695\,
            in2 => \N__22478\,
            in3 => \N__23532\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48598\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26826\,
            in1 => \N__28558\,
            in2 => \_gnd_net_\,
            in3 => \N__34608\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__23893\,
            in1 => \N__22475\,
            in2 => \N__24131\,
            in3 => \N__22463\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__22462\,
            in1 => \N__22474\,
            in2 => \N__23897\,
            in3 => \N__24130\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26827\,
            in1 => \N__28562\,
            in2 => \_gnd_net_\,
            in3 => \N__34686\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49125\,
            ce => \N__24806\,
            sr => \N__48623\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34685\,
            in1 => \N__26876\,
            in2 => \_gnd_net_\,
            in3 => \N__26894\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49125\,
            ce => \N__24806\,
            sr => \N__48623\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33922\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49119\,
            ce => 'H',
            sr => \N__48631\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33092\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33388\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33842\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33298\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33056\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33011\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33887\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48637\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23960\,
            in2 => \N__26960\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22802\,
            in2 => \N__27103\,
            in3 => \N__22784\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22781\,
            in2 => \N__27260\,
            in3 => \N__22763\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33137\,
            in2 => \N__25019\,
            in3 => \N__22724\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27202\,
            in2 => \N__22721\,
            in3 => \N__22670\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22667\,
            in2 => \N__27158\,
            in3 => \N__22628\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22625\,
            in2 => \N__27866\,
            in3 => \N__22580\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22577\,
            in2 => \N__24209\,
            in3 => \N__22541\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__49102\,
            ce => 'H',
            sr => \N__48640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33749\,
            in2 => \N__27530\,
            in3 => \N__22508\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31814\,
            in2 => \N__31868\,
            in3 => \N__22934\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22931\,
            in2 => \N__28235\,
            in3 => \N__22913\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41283\,
            in2 => \N__23123\,
            in3 => \N__22901\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22898\,
            in2 => \N__27431\,
            in3 => \N__22874\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22871\,
            in2 => \N__29915\,
            in3 => \N__22853\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31778\,
            in2 => \N__27817\,
            in3 => \N__22838\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27695\,
            in2 => \N__31796\,
            in3 => \N__22823\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__49094\,
            ce => 'H',
            sr => \N__48644\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31733\,
            in2 => \N__29840\,
            in3 => \N__22805\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27370\,
            in2 => \N__31757\,
            in3 => \N__23102\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31737\,
            in2 => \N__27638\,
            in3 => \N__23078\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35471\,
            in2 => \N__31758\,
            in3 => \N__23060\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31741\,
            in2 => \N__27749\,
            in3 => \N__23042\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27574\,
            in2 => \N__31759\,
            in3 => \N__23027\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31745\,
            in2 => \N__29984\,
            in3 => \N__23009\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29767\,
            in2 => \N__31760\,
            in3 => \N__22997\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__49085\,
            ce => 'H',
            sr => \N__48648\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31782\,
            in2 => \N__28064\,
            in3 => \N__22979\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28012\,
            in2 => \N__31797\,
            in3 => \N__22964\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31786\,
            in2 => \N__27950\,
            in3 => \N__23276\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30090\,
            in2 => \N__31798\,
            in3 => \N__23261\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31790\,
            in2 => \N__25502\,
            in3 => \N__23240\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42757\,
            in2 => \N__31799\,
            in3 => \N__23219\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31794\,
            in2 => \N__28297\,
            in3 => \N__23204\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31795\,
            in1 => \N__32033\,
            in2 => \_gnd_net_\,
            in3 => \N__23201\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49077\,
            ce => 'H',
            sr => \N__48653\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33523\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49070\,
            ce => 'H',
            sr => \N__48657\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34484\,
            in1 => \N__30403\,
            in2 => \_gnd_net_\,
            in3 => \N__30382\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30151\,
            in1 => \N__30130\,
            in2 => \_gnd_net_\,
            in3 => \N__34483\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32731\,
            in1 => \N__32707\,
            in2 => \_gnd_net_\,
            in3 => \N__34482\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__23767\,
            in1 => \N__23743\,
            in2 => \N__23300\,
            in3 => \N__23309\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__23308\,
            in1 => \N__23768\,
            in2 => \N__23747\,
            in3 => \N__23296\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28952\,
            in1 => \N__28973\,
            in2 => \_gnd_net_\,
            in3 => \N__34693\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49134\,
            ce => \N__24801\,
            sr => \N__48570\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34688\,
            in1 => \N__29012\,
            in2 => \_gnd_net_\,
            in3 => \N__29033\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49134\,
            ce => \N__24801\,
            sr => \N__48570\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29188\,
            in1 => \N__29205\,
            in2 => \_gnd_net_\,
            in3 => \N__34694\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49134\,
            ce => \N__24801\,
            sr => \N__48570\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34689\,
            in1 => \N__30274\,
            in2 => \_gnd_net_\,
            in3 => \N__30242\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49134\,
            ce => \N__24801\,
            sr => \N__48570\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28463\,
            in1 => \N__28433\,
            in2 => \_gnd_net_\,
            in3 => \N__34695\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49134\,
            ce => \N__24801\,
            sr => \N__48570\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__30147\,
            in1 => \N__30126\,
            in2 => \N__34706\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49134\,
            ce => \N__24801\,
            sr => \N__48570\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24533\,
            in2 => \N__23417\,
            in3 => \N__23533\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24527\,
            in2 => \N__23408\,
            in3 => \N__23513\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24521\,
            in2 => \N__23399\,
            in3 => \N__23720\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23390\,
            in2 => \N__23381\,
            in3 => \N__23702\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23372\,
            in2 => \N__23366\,
            in3 => \N__23684\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23663\,
            in1 => \N__23357\,
            in2 => \N__23348\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23336\,
            in2 => \N__23330\,
            in3 => \N__23642\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24425\,
            in2 => \N__23321\,
            in3 => \N__23624\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24407\,
            in2 => \N__23495\,
            in3 => \N__23606\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23486\,
            in2 => \N__24398\,
            in3 => \N__23585\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23480\,
            in2 => \N__24551\,
            in3 => \N__23867\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24557\,
            in2 => \N__23474\,
            in3 => \N__23849\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24440\,
            in2 => \N__23465\,
            in3 => \N__23831\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23810\,
            in1 => \N__24647\,
            in2 => \N__23456\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23444\,
            in2 => \N__24542\,
            in3 => \N__23792\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24329\,
            in2 => \N__24386\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23438\,
            in2 => \N__23429\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24239\,
            in2 => \N__24299\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24587\,
            in2 => \N__24641\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24974\,
            in2 => \N__24917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24902\,
            in2 => \N__24845\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23564\,
            in2 => \N__23555\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24754\,
            in2 => \N__24452\,
            in3 => \N__23543\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23540\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23537\,
            in2 => \N__24731\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24046\,
            in1 => \N__23512\,
            in2 => \_gnd_net_\,
            in3 => \N__23498\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__24050\,
            in1 => \N__23719\,
            in2 => \N__24677\,
            in3 => \N__23705\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24047\,
            in1 => \N__23701\,
            in2 => \_gnd_net_\,
            in3 => \N__23687\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24051\,
            in1 => \N__23680\,
            in2 => \_gnd_net_\,
            in3 => \N__23666\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24048\,
            in1 => \N__23659\,
            in2 => \_gnd_net_\,
            in3 => \N__23645\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24052\,
            in1 => \N__23641\,
            in2 => \_gnd_net_\,
            in3 => \N__23627\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24049\,
            in1 => \N__23623\,
            in2 => \_gnd_net_\,
            in3 => \N__23609\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48606\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24045\,
            in1 => \N__23602\,
            in2 => \_gnd_net_\,
            in3 => \N__23588\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24038\,
            in1 => \N__23581\,
            in2 => \_gnd_net_\,
            in3 => \N__23567\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24042\,
            in1 => \N__23866\,
            in2 => \_gnd_net_\,
            in3 => \N__23852\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24039\,
            in1 => \N__23848\,
            in2 => \_gnd_net_\,
            in3 => \N__23834\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24043\,
            in1 => \N__23827\,
            in2 => \_gnd_net_\,
            in3 => \N__23813\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24040\,
            in1 => \N__23809\,
            in2 => \_gnd_net_\,
            in3 => \N__23795\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24044\,
            in1 => \N__23791\,
            in2 => \_gnd_net_\,
            in3 => \N__23777\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24041\,
            in1 => \N__24370\,
            in2 => \_gnd_net_\,
            in3 => \N__23774\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49103\,
            ce => 'H',
            sr => \N__48616\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24087\,
            in1 => \N__24343\,
            in2 => \_gnd_net_\,
            in3 => \N__23771\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24098\,
            in1 => \N__23766\,
            in2 => \_gnd_net_\,
            in3 => \N__23750\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24088\,
            in1 => \N__23737\,
            in2 => \_gnd_net_\,
            in3 => \N__23723\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24099\,
            in1 => \N__24277\,
            in2 => \_gnd_net_\,
            in3 => \N__23921\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24089\,
            in1 => \N__24253\,
            in2 => \_gnd_net_\,
            in3 => \N__23918\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24100\,
            in1 => \N__24627\,
            in2 => \_gnd_net_\,
            in3 => \N__23915\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24090\,
            in1 => \N__24601\,
            in2 => \_gnd_net_\,
            in3 => \N__23912\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24101\,
            in1 => \N__24953\,
            in2 => \_gnd_net_\,
            in3 => \N__23909\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49095\,
            ce => 'H',
            sr => \N__48624\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24091\,
            in1 => \N__24933\,
            in2 => \_gnd_net_\,
            in3 => \N__23906\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24095\,
            in1 => \N__24891\,
            in2 => \_gnd_net_\,
            in3 => \N__23903\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24092\,
            in1 => \N__24870\,
            in2 => \_gnd_net_\,
            in3 => \N__23900\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24096\,
            in1 => \N__23886\,
            in2 => \_gnd_net_\,
            in3 => \N__23870\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24093\,
            in1 => \N__24121\,
            in2 => \_gnd_net_\,
            in3 => \N__24107\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24097\,
            in1 => \N__24466\,
            in2 => \_gnd_net_\,
            in3 => \N__24104\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24094\,
            in1 => \N__24490\,
            in2 => \_gnd_net_\,
            in3 => \N__23963\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33722\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49086\,
            ce => 'H',
            sr => \N__48632\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__23951\,
            in2 => \N__24158\,
            in3 => \N__23933\,
            lcout => \current_shift_inst.PI_CTRL.N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27518\,
            in1 => \N__27861\,
            in2 => \N__31864\,
            in3 => \N__24204\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__27200\,
            in1 => \N__25008\,
            in2 => \N__23939\,
            in3 => \N__27149\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23927\,
            in1 => \N__42753\,
            in2 => \N__23936\,
            in3 => \N__28233\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27685\,
            in1 => \N__41266\,
            in2 => \N__27369\,
            in3 => \N__27743\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29966\,
            in1 => \N__27630\,
            in2 => \N__35474\,
            in3 => \N__32009\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42749\,
            in2 => \_gnd_net_\,
            in3 => \N__28229\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28292\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27939\,
            in1 => \N__28004\,
            in2 => \N__28060\,
            in3 => \N__27560\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29965\,
            in1 => \N__27629\,
            in2 => \N__35473\,
            in3 => \N__28053\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30076\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27938\,
            in1 => \N__25491\,
            in2 => \N__28011\,
            in3 => \N__27559\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__24189\,
            in1 => \N__33524\,
            in2 => \N__35405\,
            in3 => \N__29486\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24188\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100010011"
        )
    port map (
            in0 => \N__32199\,
            in1 => \N__32022\,
            in2 => \N__25139\,
            in3 => \N__32381\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49065\,
            ce => 'H',
            sr => \N__48645\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__32018\,
            in1 => \N__32200\,
            in2 => \N__32398\,
            in3 => \N__25211\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49065\,
            ce => 'H',
            sr => \N__48645\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__32197\,
            in1 => \N__32020\,
            in2 => \N__25436\,
            in3 => \N__32379\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49065\,
            ce => 'H',
            sr => \N__48645\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__32019\,
            in1 => \N__32201\,
            in2 => \N__32399\,
            in3 => \N__25424\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49065\,
            ce => 'H',
            sr => \N__48645\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__32198\,
            in1 => \N__32021\,
            in2 => \N__25415\,
            in3 => \N__32380\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49065\,
            ce => 'H',
            sr => \N__48645\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27131\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100010011"
        )
    port map (
            in0 => \N__32192\,
            in1 => \N__32004\,
            in2 => \N__25175\,
            in3 => \N__32365\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49059\,
            ce => 'H',
            sr => \N__48649\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__32003\,
            in1 => \N__32193\,
            in2 => \N__32396\,
            in3 => \N__25367\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49059\,
            ce => 'H',
            sr => \N__48649\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010111"
        )
    port map (
            in0 => \N__25118\,
            in1 => \N__32366\,
            in2 => \N__32219\,
            in3 => \N__32005\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49059\,
            ce => 'H',
            sr => \N__48649\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27499\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__32028\,
            in1 => \N__32369\,
            in2 => \N__32223\,
            in3 => \N__25358\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49051\,
            ce => 'H',
            sr => \N__48654\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__32367\,
            in1 => \N__32029\,
            in2 => \N__25400\,
            in3 => \N__32211\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49051\,
            ce => 'H',
            sr => \N__48654\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__32368\,
            in1 => \N__32030\,
            in2 => \N__25388\,
            in3 => \N__32212\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49051\,
            ce => 'H',
            sr => \N__48654\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27733\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__24227\,
            in1 => \N__28154\,
            in2 => \_gnd_net_\,
            in3 => \N__28187\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49142\,
            ce => 'H',
            sr => \N__48537\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24224\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34609\,
            in1 => \N__28462\,
            in2 => \_gnd_net_\,
            in3 => \N__28422\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24226\,
            in2 => \N__28186\,
            in3 => \N__28150\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_204_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24225\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28179\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29234\,
            in1 => \N__29288\,
            in2 => \N__29184\,
            in3 => \N__28814\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26875\,
            in2 => \N__24302\,
            in3 => \N__26431\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25786\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49135\,
            ce => \N__26479\,
            sr => \N__48550\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49135\,
            ce => \N__26479\,
            sr => \N__48550\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28851\,
            in1 => \N__28815\,
            in2 => \_gnd_net_\,
            in3 => \N__34481\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29289\,
            in1 => \N__34476\,
            in2 => \_gnd_net_\,
            in3 => \N__29325\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__29235\,
            in1 => \N__29265\,
            in2 => \N__34607\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34480\,
            in1 => \N__29209\,
            in2 => \_gnd_net_\,
            in3 => \N__29177\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__24283\,
            in1 => \N__24259\,
            in2 => \N__24419\,
            in3 => \N__24434\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__24433\,
            in1 => \N__24284\,
            in2 => \N__24263\,
            in3 => \N__24415\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28895\,
            in1 => \N__28916\,
            in2 => \_gnd_net_\,
            in3 => \N__34672\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49131\,
            ce => \N__24800\,
            sr => \N__48558\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30399\,
            in1 => \N__30375\,
            in2 => \_gnd_net_\,
            in3 => \N__34673\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49131\,
            ce => \N__24800\,
            sr => \N__48558\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34768\,
            in1 => \_gnd_net_\,
            in2 => \N__34705\,
            in3 => \N__34744\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49131\,
            ce => \N__24800\,
            sr => \N__48558\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28337\,
            in1 => \N__28355\,
            in2 => \_gnd_net_\,
            in3 => \N__34674\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49131\,
            ce => \N__24800\,
            sr => \N__48558\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34668\,
            in1 => \N__32663\,
            in2 => \_gnd_net_\,
            in3 => \N__32634\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49131\,
            ce => \N__24800\,
            sr => \N__48558\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__24376\,
            in1 => \N__24352\,
            in2 => \N__24314\,
            in3 => \N__24323\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__24322\,
            in1 => \N__24377\,
            in2 => \N__24356\,
            in3 => \N__24310\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32777\,
            in1 => \N__32804\,
            in2 => \_gnd_net_\,
            in3 => \N__34679\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => \N__24802\,
            sr => \N__48571\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34675\,
            in1 => \N__32891\,
            in2 => \_gnd_net_\,
            in3 => \N__32921\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => \N__24802\,
            sr => \N__48571\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28631\,
            in1 => \N__28654\,
            in2 => \_gnd_net_\,
            in3 => \N__34678\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => \N__24802\,
            sr => \N__48571\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34676\,
            in1 => \N__28852\,
            in2 => \_gnd_net_\,
            in3 => \N__28822\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => \N__24802\,
            sr => \N__48571\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29326\,
            in1 => \N__29296\,
            in2 => \_gnd_net_\,
            in3 => \N__34680\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => \N__24802\,
            sr => \N__48571\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34677\,
            in1 => \N__29236\,
            in2 => \_gnd_net_\,
            in3 => \N__29266\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => \N__24802\,
            sr => \N__48571\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__24474\,
            in1 => \N__24660\,
            in2 => \N__24503\,
            in3 => \N__24514\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__24513\,
            in1 => \N__24501\,
            in2 => \N__24664\,
            in3 => \N__24475\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28493\,
            in1 => \N__28792\,
            in2 => \_gnd_net_\,
            in3 => \N__34616\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49120\,
            ce => \N__24803\,
            sr => \N__48581\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__24515\,
            in1 => \N__24502\,
            in2 => \N__24665\,
            in3 => \N__24476\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28687\,
            in1 => \N__34614\,
            in2 => \_gnd_net_\,
            in3 => \N__28674\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28675\,
            in1 => \_gnd_net_\,
            in2 => \N__24443\,
            in3 => \N__34622\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49120\,
            ce => \N__24803\,
            sr => \N__48581\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34623\,
            in1 => \N__28769\,
            in2 => \_gnd_net_\,
            in3 => \N__28744\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49120\,
            ce => \N__24803\,
            sr => \N__48581\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34615\,
            in1 => \N__32842\,
            in2 => \_gnd_net_\,
            in3 => \N__32867\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49120\,
            ce => \N__24803\,
            sr => \N__48581\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__24628\,
            in1 => \N__24607\,
            in2 => \N__24572\,
            in3 => \N__24581\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__24580\,
            in1 => \N__24629\,
            in2 => \N__24611\,
            in3 => \N__24568\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32735\,
            in1 => \N__32699\,
            in2 => \_gnd_net_\,
            in3 => \N__34667\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49112\,
            ce => \N__24804\,
            sr => \N__48588\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34664\,
            in1 => \_gnd_net_\,
            in2 => \N__30197\,
            in3 => \N__30218\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49112\,
            ce => \N__24804\,
            sr => \N__48588\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28606\,
            in1 => \N__34662\,
            in2 => \_gnd_net_\,
            in3 => \N__28573\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34663\,
            in1 => \_gnd_net_\,
            in2 => \N__24560\,
            in3 => \N__28607\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49112\,
            ce => \N__24804\,
            sr => \N__48588\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28385\,
            in1 => \N__34666\,
            in2 => \_gnd_net_\,
            in3 => \N__28406\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49112\,
            ce => \N__24804\,
            sr => \N__48588\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34665\,
            in1 => \N__29073\,
            in2 => \_gnd_net_\,
            in3 => \N__29093\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49112\,
            ce => \N__24804\,
            sr => \N__48588\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__27035\,
            in1 => \N__35743\,
            in2 => \N__27053\,
            in3 => \N__26987\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__26678\,
            in1 => \N__24718\,
            in2 => \N__24779\,
            in3 => \N__34841\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49104\,
            ce => 'H',
            sr => \N__48599\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__26785\,
            in1 => \N__24775\,
            in2 => \_gnd_net_\,
            in3 => \N__24713\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__24776\,
            in1 => \N__26758\,
            in2 => \N__26744\,
            in3 => \N__26787\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49104\,
            ce => 'H',
            sr => \N__48599\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__26786\,
            in1 => \N__24767\,
            in2 => \N__24758\,
            in3 => \N__24740\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24734\,
            in3 => \N__26728\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24714\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49104\,
            ce => 'H',
            sr => \N__48599\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26729\,
            in2 => \_gnd_net_\,
            in3 => \N__24688\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__24951\,
            in1 => \N__24934\,
            in2 => \N__24818\,
            in3 => \N__24965\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__24964\,
            in1 => \N__24952\,
            in2 => \N__24938\,
            in3 => \N__24814\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29446\,
            in1 => \N__29416\,
            in2 => \_gnd_net_\,
            in3 => \N__34696\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34698\,
            in1 => \_gnd_net_\,
            in2 => \N__24905\,
            in3 => \N__29447\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49096\,
            ce => \N__24805\,
            sr => \N__48607\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__24853\,
            in1 => \N__24893\,
            in2 => \N__24875\,
            in3 => \N__24826\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__24892\,
            in1 => \N__24871\,
            in2 => \N__24830\,
            in3 => \N__24854\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26432\,
            in1 => \N__26444\,
            in2 => \_gnd_net_\,
            in3 => \N__34699\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49096\,
            ce => \N__24805\,
            sr => \N__48607\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34697\,
            in1 => \N__29141\,
            in2 => \_gnd_net_\,
            in3 => \N__29156\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49096\,
            ce => \N__24805\,
            sr => \N__48607\
        );

    \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__24993\,
            in1 => \N__33838\,
            in2 => \N__35380\,
            in3 => \N__29534\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24992\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010111111111"
        )
    port map (
            in0 => \N__32158\,
            in1 => \_gnd_net_\,
            in2 => \N__32395\,
            in3 => \N__25031\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49087\,
            ce => 'H',
            sr => \N__48617\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__32013\,
            in1 => \N__32350\,
            in2 => \N__32202\,
            in3 => \N__25100\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49087\,
            ce => 'H',
            sr => \N__48617\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011111110"
        )
    port map (
            in0 => \N__32156\,
            in1 => \N__32016\,
            in2 => \N__32393\,
            in3 => \N__25079\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49087\,
            ce => 'H',
            sr => \N__48617\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__32014\,
            in1 => \N__32351\,
            in2 => \N__32203\,
            in3 => \N__25349\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49087\,
            ce => 'H',
            sr => \N__48617\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011111110"
        )
    port map (
            in0 => \N__32157\,
            in1 => \N__32017\,
            in2 => \N__32394\,
            in3 => \N__25337\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49087\,
            ce => 'H',
            sr => \N__48617\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__32015\,
            in1 => \N__32352\,
            in2 => \N__32204\,
            in3 => \N__25313\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49087\,
            ce => 'H',
            sr => \N__48617\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27193\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__32132\,
            in1 => \N__32027\,
            in2 => \N__25196\,
            in3 => \N__32328\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49078\,
            ce => 'H',
            sr => \N__48625\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__32023\,
            in1 => \N__32133\,
            in2 => \N__32382\,
            in3 => \N__25301\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49078\,
            ce => 'H',
            sr => \N__48625\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__32130\,
            in1 => \N__32025\,
            in2 => \N__25280\,
            in3 => \N__32326\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49078\,
            ce => 'H',
            sr => \N__48625\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__32024\,
            in1 => \N__32134\,
            in2 => \N__32383\,
            in3 => \N__25250\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49078\,
            ce => 'H',
            sr => \N__48625\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__32131\,
            in1 => \N__32026\,
            in2 => \N__25238\,
            in3 => \N__32327\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49078\,
            ce => 'H',
            sr => \N__48625\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27271\,
            in2 => \N__27275\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26930\,
            in2 => \N__26918\,
            in3 => \N__25064\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27281\,
            in2 => \N__27065\,
            in3 => \N__25061\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27227\,
            in2 => \N__27290\,
            in3 => \N__25058\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25055\,
            in2 => \N__25046\,
            in3 => \N__25022\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25202\,
            in2 => \N__27167\,
            in3 => \N__25187\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25184\,
            in2 => \N__27113\,
            in3 => \N__25160\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27959\,
            in2 => \N__27887\,
            in3 => \N__25157\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25154\,
            in2 => \N__25148\,
            in3 => \N__25130\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25127\,
            in2 => \N__27476\,
            in3 => \N__25109\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27644\,
            in2 => \N__27221\,
            in3 => \N__25106\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28070\,
            in2 => \N__27452\,
            in3 => \N__25103\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41225\,
            in2 => \N__27443\,
            in3 => \N__25091\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25088\,
            in2 => \N__27380\,
            in3 => \N__25067\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27467\,
            in2 => \N__29867\,
            in3 => \N__25340\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27767\,
            in2 => \N__27461\,
            in3 => \N__25328\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25325\,
            in2 => \N__27653\,
            in3 => \N__25304\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29777\,
            in2 => \N__27584\,
            in3 => \N__25292\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25289\,
            in2 => \N__27323\,
            in3 => \N__25268\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25265\,
            in2 => \N__27593\,
            in3 => \N__25241\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35420\,
            in2 => \N__27308\,
            in3 => \N__25226\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25223\,
            in2 => \N__27704\,
            in3 => \N__25205\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27536\,
            in2 => \N__27761\,
            in3 => \N__25427\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29945\,
            in2 => \N__27899\,
            in3 => \N__25418\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29852\,
            in2 => \N__29708\,
            in3 => \N__25406\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25523\,
            in2 => \N__28022\,
            in3 => \N__25403\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25511\,
            in2 => \N__27968\,
            in3 => \N__25391\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25517\,
            in2 => \N__27908\,
            in3 => \N__25379\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25376\,
            in2 => \N__30041\,
            in3 => \N__25361\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25460\,
            in2 => \N__30316\,
            in3 => \N__25352\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30312\,
            in2 => \N__42710\,
            in3 => \N__25541\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25538\,
            in2 => \N__30317\,
            in3 => \N__25529\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35402\,
            in1 => \N__31922\,
            in2 => \_gnd_net_\,
            in3 => \N__25526\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28043\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27931\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27994\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25487\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__31992\,
            in1 => \N__32397\,
            in2 => \N__32224\,
            in3 => \N__25454\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49036\,
            ce => 'H',
            sr => \N__48655\
        );

    \phase_controller_inst2.S2_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26996\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49036\,
            ce => 'H',
            sr => \N__48655\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25942\,
            in1 => \N__25776\,
            in2 => \_gnd_net_\,
            in3 => \N__25568\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25938\,
            in1 => \N__25749\,
            in2 => \_gnd_net_\,
            in3 => \N__25565\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25943\,
            in1 => \N__25726\,
            in2 => \_gnd_net_\,
            in3 => \N__25562\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25939\,
            in1 => \N__25698\,
            in2 => \_gnd_net_\,
            in3 => \N__25559\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25944\,
            in1 => \N__25668\,
            in2 => \_gnd_net_\,
            in3 => \N__25556\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25940\,
            in1 => \N__25641\,
            in2 => \_gnd_net_\,
            in3 => \N__25553\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25945\,
            in1 => \N__26161\,
            in2 => \_gnd_net_\,
            in3 => \N__25550\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25941\,
            in1 => \N__26137\,
            in2 => \_gnd_net_\,
            in3 => \N__25547\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__49143\,
            ce => \N__25829\,
            sr => \N__48527\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25927\,
            in1 => \N__26106\,
            in2 => \_gnd_net_\,
            in3 => \N__25544\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25931\,
            in1 => \N__26079\,
            in2 => \_gnd_net_\,
            in3 => \N__25595\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25924\,
            in1 => \N__26050\,
            in2 => \_gnd_net_\,
            in3 => \N__25592\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25928\,
            in1 => \N__26022\,
            in2 => \_gnd_net_\,
            in3 => \N__25589\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25925\,
            in1 => \N__25995\,
            in2 => \_gnd_net_\,
            in3 => \N__25586\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25929\,
            in1 => \N__25974\,
            in2 => \_gnd_net_\,
            in3 => \N__25583\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25926\,
            in1 => \N__26392\,
            in2 => \_gnd_net_\,
            in3 => \N__25580\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25930\,
            in1 => \N__26367\,
            in2 => \_gnd_net_\,
            in3 => \N__25577\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__49139\,
            ce => \N__25818\,
            sr => \N__48531\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25920\,
            in1 => \N__26334\,
            in2 => \_gnd_net_\,
            in3 => \N__25574\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25946\,
            in1 => \N__26307\,
            in2 => \_gnd_net_\,
            in3 => \N__25571\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25921\,
            in1 => \N__26283\,
            in2 => \_gnd_net_\,
            in3 => \N__25622\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25947\,
            in1 => \N__26262\,
            in2 => \_gnd_net_\,
            in3 => \N__25619\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25922\,
            in1 => \N__26235\,
            in2 => \_gnd_net_\,
            in3 => \N__25616\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25948\,
            in1 => \N__26208\,
            in2 => \_gnd_net_\,
            in3 => \N__25613\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25923\,
            in1 => \N__26182\,
            in2 => \_gnd_net_\,
            in3 => \N__25610\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25949\,
            in1 => \N__26658\,
            in2 => \_gnd_net_\,
            in3 => \N__25607\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__49136\,
            ce => \N__25809\,
            sr => \N__48538\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25932\,
            in1 => \N__26625\,
            in2 => \_gnd_net_\,
            in3 => \N__25604\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__49132\,
            ce => \N__25825\,
            sr => \N__48544\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25936\,
            in1 => \N__26601\,
            in2 => \_gnd_net_\,
            in3 => \N__25601\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__49132\,
            ce => \N__25825\,
            sr => \N__48544\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25933\,
            in1 => \N__26577\,
            in2 => \_gnd_net_\,
            in3 => \N__25598\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__49132\,
            ce => \N__25825\,
            sr => \N__48544\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25937\,
            in1 => \N__26517\,
            in2 => \_gnd_net_\,
            in3 => \N__25955\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__49132\,
            ce => \N__25825\,
            sr => \N__48544\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25934\,
            in1 => \N__26557\,
            in2 => \_gnd_net_\,
            in3 => \N__25952\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__49132\,
            ce => \N__25825\,
            sr => \N__48544\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26536\,
            in1 => \N__25935\,
            in2 => \_gnd_net_\,
            in3 => \N__25832\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49132\,
            ce => \N__25825\,
            sr => \N__48544\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25732\,
            in2 => \N__25787\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25756\,
            in2 => \N__25709\,
            in3 => \N__25736\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25733\,
            in2 => \N__25675\,
            in3 => \N__25712\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25708\,
            in2 => \N__25648\,
            in3 => \N__25679\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26167\,
            in2 => \N__25676\,
            in3 => \N__25652\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26143\,
            in2 => \N__25649\,
            in3 => \N__25625\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26168\,
            in2 => \N__26119\,
            in3 => \N__26147\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26144\,
            in2 => \N__26086\,
            in3 => \N__26123\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49127\,
            ce => \N__26490\,
            sr => \N__48551\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26056\,
            in2 => \N__26120\,
            in3 => \N__26090\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26029\,
            in2 => \N__26087\,
            in3 => \N__26060\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26057\,
            in2 => \N__26002\,
            in3 => \N__26036\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25975\,
            in2 => \N__26033\,
            in3 => \N__26006\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26398\,
            in2 => \N__26003\,
            in3 => \N__25979\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25976\,
            in2 => \N__26374\,
            in3 => \N__25958\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26399\,
            in2 => \N__26347\,
            in3 => \N__26378\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26308\,
            in2 => \N__26375\,
            in3 => \N__26351\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49121\,
            ce => \N__26483\,
            sr => \N__48559\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26284\,
            in2 => \N__26348\,
            in3 => \N__26318\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26263\,
            in2 => \N__26315\,
            in3 => \N__26288\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26285\,
            in2 => \N__26242\,
            in3 => \N__26267\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26264\,
            in2 => \N__26215\,
            in3 => \N__26246\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26188\,
            in2 => \N__26243\,
            in3 => \N__26219\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26665\,
            in2 => \N__26216\,
            in3 => \N__26192\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26189\,
            in2 => \N__26638\,
            in3 => \N__26672\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26602\,
            in2 => \N__26669\,
            in3 => \N__26642\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49113\,
            ce => \N__26491\,
            sr => \N__48572\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26578\,
            in2 => \N__26639\,
            in3 => \N__26609\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49105\,
            ce => \N__26492\,
            sr => \N__48582\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26518\,
            in2 => \N__26606\,
            in3 => \N__26582\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49105\,
            ce => \N__26492\,
            sr => \N__48582\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26579\,
            in2 => \N__26561\,
            in3 => \N__26543\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49105\,
            ce => \N__26492\,
            sr => \N__48582\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26540\,
            in2 => \N__26522\,
            in3 => \N__26498\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49105\,
            ce => \N__26492\,
            sr => \N__48582\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26495\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49105\,
            ce => \N__26492\,
            sr => \N__48582\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26423\,
            in1 => \N__26443\,
            in2 => \_gnd_net_\,
            in3 => \N__34701\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__34702\,
            in1 => \N__26424\,
            in2 => \N__26402\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49097\,
            ce => \N__34242\,
            sr => \N__48589\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26864\,
            in1 => \N__26890\,
            in2 => \_gnd_net_\,
            in3 => \N__34700\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34703\,
            in1 => \_gnd_net_\,
            in2 => \N__26879\,
            in3 => \N__26865\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49097\,
            ce => \N__34242\,
            sr => \N__48589\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__26803\,
            in1 => \N__30931\,
            in2 => \N__26843\,
            in3 => \N__30538\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__30932\,
            in1 => \N__26804\,
            in2 => \N__30539\,
            in3 => \N__26842\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26831\,
            in1 => \N__28547\,
            in2 => \_gnd_net_\,
            in3 => \N__34704\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49097\,
            ce => \N__34242\,
            sr => \N__48589\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__29405\,
            in1 => \N__30563\,
            in2 => \N__30596\,
            in3 => \N__29393\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__26988\,
            in1 => \N__27033\,
            in2 => \N__26693\,
            in3 => \N__26705\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49088\,
            ce => 'H',
            sr => \N__48600\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010101010"
        )
    port map (
            in0 => \N__26704\,
            in1 => \N__26791\,
            in2 => \N__26765\,
            in3 => \N__26736\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49088\,
            ce => 'H',
            sr => \N__48600\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26703\,
            in2 => \_gnd_net_\,
            in3 => \N__26689\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__31649\,
            in1 => \N__31681\,
            in2 => \N__27056\,
            in3 => \N__33659\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49088\,
            ce => 'H',
            sr => \N__48600\
        );

    \phase_controller_inst2.state_2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__27049\,
            in1 => \N__31680\,
            in2 => \N__35744\,
            in3 => \N__31650\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49088\,
            ce => 'H',
            sr => \N__48600\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27048\,
            in2 => \_gnd_net_\,
            in3 => \N__35739\,
            lcout => \phase_controller_inst2.state_RNIG7JFZ0Z_2\,
            ltout => \phase_controller_inst2.state_RNIG7JFZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__27034\,
            in1 => \_gnd_net_\,
            in2 => \N__26999\,
            in3 => \N__26989\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49088\,
            ce => 'H',
            sr => \N__48600\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__32390\,
            in1 => \N__32154\,
            in2 => \_gnd_net_\,
            in3 => \N__26969\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49079\,
            ce => 'H',
            sr => \N__48608\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33006\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26941\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => \current_shift_inst.PI_CTRL.integrator_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35292\,
            in1 => \N__33007\,
            in2 => \N__26921\,
            in3 => \N__29351\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__32391\,
            in1 => \N__32155\,
            in2 => \_gnd_net_\,
            in3 => \N__26903\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49079\,
            ce => 'H',
            sr => \N__48608\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__32153\,
            in1 => \N__32392\,
            in2 => \_gnd_net_\,
            in3 => \N__27299\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49079\,
            ce => 'H',
            sr => \N__48608\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35336\,
            in1 => \N__27241\,
            in2 => \N__33886\,
            in3 => \N__29543\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27083\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35339\,
            in1 => \N__31857\,
            in2 => \N__33299\,
            in3 => \N__29456\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__27201\,
            in1 => \N__35337\,
            in2 => \N__29522\,
            in3 => \N__33964\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35338\,
            in1 => \N__27157\,
            in2 => \N__33482\,
            in3 => \N__29510\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__33923\,
            in1 => \N__35335\,
            in2 => \N__29342\,
            in3 => \N__27084\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__33188\,
            in1 => \N__27528\,
            in2 => \N__35397\,
            in3 => \N__29465\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33187\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__29909\,
            in1 => \N__35354\,
            in2 => \N__33416\,
            in3 => \N__29603\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__27818\,
            in1 => \N__35368\,
            in2 => \N__31469\,
            in3 => \N__29594\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__28234\,
            in1 => \N__29630\,
            in2 => \N__35398\,
            in3 => \N__33347\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__41276\,
            in1 => \N__33323\,
            in2 => \N__35395\,
            in3 => \N__29621\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__27409\,
            in1 => \N__33440\,
            in2 => \N__35399\,
            in3 => \N__29612\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__27352\,
            in1 => \N__35129\,
            in2 => \N__35396\,
            in3 => \N__29561\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__35461\,
            in1 => \N__30024\,
            in2 => \N__35384\,
            in3 => \N__29696\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27808\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__31418\,
            in2 => \N__35383\,
            in3 => \N__29678\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__27748\,
            in1 => \N__35330\,
            in2 => \N__32435\,
            in3 => \N__29687\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__27694\,
            in1 => \N__32459\,
            in2 => \N__35381\,
            in3 => \N__29585\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__27634\,
            in1 => \N__32483\,
            in2 => \N__35382\,
            in3 => \N__29552\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__31493\,
            in1 => \N__29839\,
            in2 => \N__29576\,
            in3 => \N__35320\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27567\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28205\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__31445\,
            in1 => \N__28052\,
            in2 => \N__35401\,
            in3 => \N__29657\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__28013\,
            in1 => \N__35375\,
            in2 => \N__29936\,
            in3 => \N__29648\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__27949\,
            in1 => \N__35376\,
            in2 => \N__30005\,
            in3 => \N__29639\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__32507\,
            in1 => \N__29977\,
            in2 => \N__35400\,
            in3 => \N__29669\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__27854\,
            in1 => \N__33389\,
            in2 => \N__35403\,
            in3 => \N__29501\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111011101"
        )
    port map (
            in0 => \N__31947\,
            in1 => \N__32389\,
            in2 => \N__32215\,
            in3 => \N__27875\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49046\,
            ce => 'H',
            sr => \N__48641\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__31945\,
            in1 => \N__32387\,
            in2 => \N__32213\,
            in3 => \N__27824\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49046\,
            ce => 'H',
            sr => \N__48641\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__32386\,
            in1 => \N__31949\,
            in2 => \N__28319\,
            in3 => \N__32188\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49046\,
            ce => 'H',
            sr => \N__48641\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__31946\,
            in1 => \N__32388\,
            in2 => \N__32214\,
            in3 => \N__28307\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49046\,
            ce => 'H',
            sr => \N__48641\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__32385\,
            in1 => \N__31948\,
            in2 => \N__28253\,
            in3 => \N__32187\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49046\,
            ce => 'H',
            sr => \N__48641\
        );

    \delay_measurement_inst.stop_timer_tr_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28135\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28118\,
            ce => 'H',
            sr => \N__48646\
        );

    \delay_measurement_inst.start_timer_tr_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28134\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28118\,
            ce => 'H',
            sr => \N__48646\
        );

    \phase_controller_inst2.S1_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31654\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49017\,
            ce => 'H',
            sr => \N__48658\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30238\,
            in1 => \N__30273\,
            in2 => \_gnd_net_\,
            in3 => \N__34532\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30368\,
            in2 => \_gnd_net_\,
            in3 => \N__30113\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28454\,
            in1 => \N__30263\,
            in2 => \N__28478\,
            in3 => \N__28361\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__28475\,
            in1 => \N__28748\,
            in2 => \N__28466\,
            in3 => \N__28520\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28455\,
            in1 => \_gnd_net_\,
            in2 => \N__28436\,
            in3 => \N__28429\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49122\,
            ce => \N__34199\,
            sr => \N__48532\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34468\,
            in1 => \N__28381\,
            in2 => \_gnd_net_\,
            in3 => \N__28399\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28380\,
            in2 => \N__28388\,
            in3 => \N__34472\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49114\,
            ce => \N__34183\,
            sr => \N__48539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28379\,
            in1 => \N__32630\,
            in2 => \N__28605\,
            in3 => \N__28334\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28335\,
            in1 => \N__28351\,
            in2 => \_gnd_net_\,
            in3 => \N__34469\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34470\,
            in1 => \_gnd_net_\,
            in2 => \N__28340\,
            in3 => \N__28336\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49114\,
            ce => \N__34183\,
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28604\,
            in1 => \N__34471\,
            in2 => \_gnd_net_\,
            in3 => \N__28580\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49114\,
            ce => \N__34183\,
            sr => \N__48539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28793\,
            in1 => \N__29433\,
            in2 => \N__28557\,
            in3 => \N__29124\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28499\,
            in1 => \N__28505\,
            in2 => \N__28523\,
            in3 => \N__28511\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28649\,
            in1 => \N__32838\,
            in2 => \N__32805\,
            in3 => \N__28673\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29003\,
            in1 => \N__28938\,
            in2 => \N__32922\,
            in3 => \N__28884\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30180\,
            in1 => \N__29067\,
            in2 => \N__32700\,
            in3 => \N__34724\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28629\,
            in1 => \N__28650\,
            in2 => \_gnd_net_\,
            in3 => \N__34598\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100001010"
        )
    port map (
            in0 => \N__30880\,
            in1 => \N__30906\,
            in2 => \N__28720\,
            in3 => \N__28702\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28790\,
            in1 => \N__34511\,
            in2 => \_gnd_net_\,
            in3 => \N__28489\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34513\,
            in1 => \_gnd_net_\,
            in2 => \N__28796\,
            in3 => \N__28791\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49098\,
            ce => \N__34259\,
            sr => \N__48552\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28742\,
            in1 => \_gnd_net_\,
            in2 => \N__28768\,
            in3 => \N__34512\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => \elapsed_time_ns_1_RNI0CQBB_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34514\,
            in1 => \_gnd_net_\,
            in2 => \N__28751\,
            in3 => \N__28743\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49098\,
            ce => \N__34259\,
            sr => \N__48552\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28703\,
            in1 => \N__28719\,
            in2 => \N__30911\,
            in3 => \N__30881\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__30879\,
            in1 => \N__30907\,
            in2 => \N__28721\,
            in3 => \N__28701\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28691\,
            in1 => \N__34515\,
            in2 => \_gnd_net_\,
            in3 => \N__28676\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49098\,
            ce => \N__34259\,
            sr => \N__48552\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__30475\,
            in1 => \N__30492\,
            in2 => \N__28985\,
            in3 => \N__28925\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28655\,
            in1 => \N__28630\,
            in2 => \_gnd_net_\,
            in3 => \N__34591\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49090\,
            ce => \N__34250\,
            sr => \N__48563\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28924\,
            in1 => \N__30474\,
            in2 => \N__30497\,
            in3 => \N__28981\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29004\,
            in1 => \N__29026\,
            in2 => \_gnd_net_\,
            in3 => \N__34588\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34590\,
            in1 => \_gnd_net_\,
            in2 => \N__29015\,
            in3 => \N__29005\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49090\,
            ce => \N__34250\,
            sr => \N__48563\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28947\,
            in1 => \N__28966\,
            in2 => \_gnd_net_\,
            in3 => \N__34587\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34589\,
            in1 => \_gnd_net_\,
            in2 => \N__28955\,
            in3 => \N__28948\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49090\,
            ce => \N__34250\,
            sr => \N__48563\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__30456\,
            in1 => \N__28868\,
            in2 => \N__34274\,
            in3 => \N__30702\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28893\,
            in1 => \N__28909\,
            in2 => \_gnd_net_\,
            in3 => \N__34592\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34594\,
            in1 => \_gnd_net_\,
            in2 => \N__28898\,
            in3 => \N__28894\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49081\,
            ce => \N__34244\,
            sr => \N__48573\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__28867\,
            in1 => \N__34273\,
            in2 => \N__30707\,
            in3 => \N__30457\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34593\,
            in1 => \N__28859\,
            in2 => \_gnd_net_\,
            in3 => \N__28829\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49081\,
            ce => \N__34244\,
            sr => \N__48573\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29330\,
            in1 => \N__29303\,
            in2 => \_gnd_net_\,
            in3 => \N__34596\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49081\,
            ce => \N__34244\,
            sr => \N__48573\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34595\,
            in1 => \N__29270\,
            in2 => \_gnd_net_\,
            in3 => \N__29243\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49081\,
            ce => \N__34244\,
            sr => \N__48573\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29216\,
            in1 => \N__29189\,
            in2 => \_gnd_net_\,
            in3 => \N__34597\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49081\,
            ce => \N__34244\,
            sr => \N__48573\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__29044\,
            in1 => \N__30615\,
            in2 => \N__29105\,
            in3 => \N__30638\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100110001"
        )
    port map (
            in0 => \N__30637\,
            in1 => \N__30616\,
            in2 => \N__29048\,
            in3 => \N__29101\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34602\,
            in1 => \N__29139\,
            in2 => \_gnd_net_\,
            in3 => \N__29152\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29140\,
            in1 => \_gnd_net_\,
            in2 => \N__29108\,
            in3 => \N__34605\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49071\,
            ce => \N__34245\,
            sr => \N__48583\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29074\,
            in1 => \_gnd_net_\,
            in2 => \N__34684\,
            in3 => \N__29086\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29075\,
            in2 => \N__29051\,
            in3 => \N__34604\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49071\,
            ce => \N__34245\,
            sr => \N__48583\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34603\,
            in1 => \N__29445\,
            in2 => \_gnd_net_\,
            in3 => \N__29420\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49071\,
            ce => \N__34245\,
            sr => \N__48583\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__29404\,
            in1 => \N__30558\,
            in2 => \N__30592\,
            in3 => \N__29392\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29381\,
            in2 => \_gnd_net_\,
            in3 => \N__33715\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29375\,
            in2 => \_gnd_net_\,
            in3 => \N__33088\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29369\,
            in2 => \_gnd_net_\,
            in3 => \N__33052\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29363\,
            in2 => \_gnd_net_\,
            in3 => \N__33155\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29357\,
            in2 => \_gnd_net_\,
            in3 => \N__29345\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33896\,
            in2 => \_gnd_net_\,
            in3 => \N__29333\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33851\,
            in2 => \_gnd_net_\,
            in3 => \N__29537\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33812\,
            in2 => \_gnd_net_\,
            in3 => \N__29525\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33935\,
            in2 => \_gnd_net_\,
            in3 => \N__29513\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33449\,
            in2 => \_gnd_net_\,
            in3 => \N__29504\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33356\,
            in2 => \_gnd_net_\,
            in3 => \N__29489\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33491\,
            in2 => \_gnd_net_\,
            in3 => \N__29474\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29471\,
            in2 => \_gnd_net_\,
            in3 => \N__29459\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33266\,
            in2 => \_gnd_net_\,
            in3 => \N__29450\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33343\,
            in2 => \_gnd_net_\,
            in3 => \N__29624\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33319\,
            in2 => \_gnd_net_\,
            in3 => \N__29615\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33439\,
            in2 => \_gnd_net_\,
            in3 => \N__29606\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33412\,
            in2 => \_gnd_net_\,
            in3 => \N__29597\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31461\,
            in2 => \_gnd_net_\,
            in3 => \N__29588\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32451\,
            in2 => \_gnd_net_\,
            in3 => \N__29579\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31485\,
            in2 => \_gnd_net_\,
            in3 => \N__29564\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35128\,
            in2 => \_gnd_net_\,
            in3 => \N__29555\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32475\,
            in2 => \_gnd_net_\,
            in3 => \N__29546\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30026\,
            in2 => \_gnd_net_\,
            in3 => \N__29690\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32424\,
            in2 => \_gnd_net_\,
            in3 => \N__29681\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31410\,
            in2 => \_gnd_net_\,
            in3 => \N__29672\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32499\,
            in2 => \_gnd_net_\,
            in3 => \N__29663\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33637\,
            in2 => \_gnd_net_\,
            in3 => \N__29660\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31441\,
            in3 => \N__29651\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29931\,
            in2 => \_gnd_net_\,
            in3 => \N__29642\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30000\,
            in2 => \_gnd_net_\,
            in3 => \N__29633\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__30094\,
            in1 => \N__35358\,
            in2 => \_gnd_net_\,
            in3 => \N__30044\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30025\,
            in2 => \_gnd_net_\,
            in3 => \N__35331\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35333\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29976\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35332\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29908\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29755\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29824\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__33641\,
            in1 => \N__29768\,
            in2 => \N__35404\,
            in3 => \N__29717\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35391\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30284\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30278\,
            in1 => \N__30234\,
            in2 => \_gnd_net_\,
            in3 => \N__34606\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49129\,
            ce => \N__34251\,
            sr => \N__48521\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__30659\,
            in1 => \N__30682\,
            in2 => \N__30164\,
            in3 => \N__32672\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__32671\,
            in1 => \N__30658\,
            in2 => \N__30686\,
            in3 => \N__30160\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30195\,
            in1 => \N__34575\,
            in2 => \_gnd_net_\,
            in3 => \N__30211\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34576\,
            in1 => \_gnd_net_\,
            in2 => \N__30200\,
            in3 => \N__30196\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49115\,
            ce => \N__34243\,
            sr => \N__48528\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30152\,
            in1 => \N__30131\,
            in2 => \_gnd_net_\,
            in3 => \N__34578\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49115\,
            ce => \N__34243\,
            sr => \N__48528\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34577\,
            in1 => \N__30404\,
            in2 => \_gnd_net_\,
            in3 => \N__30383\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49115\,
            ce => \N__34243\,
            sr => \N__48528\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35099\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49107\,
            ce => 'H',
            sr => \N__48533\
        );

    \phase_controller_inst1.stoper_tr.running_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000111010"
        )
    port map (
            in0 => \N__30338\,
            in1 => \N__34962\,
            in2 => \N__34941\,
            in3 => \N__35003\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49107\,
            ce => 'H',
            sr => \N__48533\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__34961\,
            in1 => \N__30350\,
            in2 => \N__31531\,
            in3 => \N__31511\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30341\,
            in3 => \N__34925\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__34960\,
            in1 => \N__30337\,
            in2 => \_gnd_net_\,
            in3 => \N__35098\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30329\,
            in3 => \N__30856\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30326\,
            in2 => \N__30839\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34175\,
            in1 => \N__30793\,
            in2 => \_gnd_net_\,
            in3 => \N__30320\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__34252\,
            in1 => \N__30766\,
            in2 => \N__30440\,
            in3 => \N__30431\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34176\,
            in1 => \N__30727\,
            in2 => \_gnd_net_\,
            in3 => \N__30428\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34253\,
            in1 => \N__31186\,
            in2 => \_gnd_net_\,
            in3 => \N__30425\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34177\,
            in1 => \N__31147\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34254\,
            in1 => \N__31096\,
            in2 => \_gnd_net_\,
            in3 => \N__30419\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34178\,
            in1 => \N__31057\,
            in2 => \_gnd_net_\,
            in3 => \N__30416\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49099\,
            ce => 'H',
            sr => \N__48540\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34182\,
            in1 => \N__31018\,
            in2 => \_gnd_net_\,
            in3 => \N__30413\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34163\,
            in1 => \N__30994\,
            in2 => \_gnd_net_\,
            in3 => \N__30410\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34179\,
            in1 => \N__30955\,
            in2 => \_gnd_net_\,
            in3 => \N__30407\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34164\,
            in1 => \N__31378\,
            in2 => \_gnd_net_\,
            in3 => \N__30515\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34180\,
            in1 => \N__31357\,
            in2 => \_gnd_net_\,
            in3 => \N__30512\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34165\,
            in1 => \N__31318\,
            in2 => \_gnd_net_\,
            in3 => \N__30509\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34181\,
            in1 => \N__31294\,
            in2 => \_gnd_net_\,
            in3 => \N__30506\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34166\,
            in1 => \N__32564\,
            in2 => \_gnd_net_\,
            in3 => \N__30503\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49091\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34246\,
            in1 => \N__32584\,
            in2 => \_gnd_net_\,
            in3 => \N__30500\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34189\,
            in1 => \N__30496\,
            in2 => \_gnd_net_\,
            in3 => \N__30479\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34247\,
            in1 => \N__30476\,
            in2 => \_gnd_net_\,
            in3 => \N__30461\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34190\,
            in1 => \N__30458\,
            in2 => \_gnd_net_\,
            in3 => \N__30443\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34248\,
            in1 => \N__30706\,
            in2 => \_gnd_net_\,
            in3 => \N__30689\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34191\,
            in1 => \N__30676\,
            in2 => \_gnd_net_\,
            in3 => \N__30662\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34249\,
            in1 => \N__30657\,
            in2 => \_gnd_net_\,
            in3 => \N__30641\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__30636\,
            in2 => \_gnd_net_\,
            in3 => \N__30620\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49082\,
            ce => 'H',
            sr => \N__48553\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34200\,
            in1 => \N__30617\,
            in2 => \_gnd_net_\,
            in3 => \N__30599\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34205\,
            in1 => \N__30588\,
            in2 => \_gnd_net_\,
            in3 => \N__30566\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34201\,
            in1 => \N__30562\,
            in2 => \_gnd_net_\,
            in3 => \N__30542\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34206\,
            in1 => \N__30534\,
            in2 => \_gnd_net_\,
            in3 => \N__30518\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34202\,
            in1 => \N__30930\,
            in2 => \_gnd_net_\,
            in3 => \N__30914\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34207\,
            in1 => \N__30905\,
            in2 => \_gnd_net_\,
            in3 => \N__30887\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34203\,
            in1 => \N__30878\,
            in2 => \_gnd_net_\,
            in3 => \N__30884\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__34943\,
            in1 => \N__30860\,
            in2 => \N__30835\,
            in3 => \N__34204\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49072\,
            ce => 'H',
            sr => \N__48564\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30845\,
            in2 => \N__30809\,
            in3 => \N__30825\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30800\,
            in2 => \N__30779\,
            in3 => \N__30794\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30770\,
            in1 => \N__30752\,
            in2 => \N__30746\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30713\,
            in2 => \N__30737\,
            in3 => \N__30728\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31187\,
            in1 => \N__31172\,
            in2 => \N__31157\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31148\,
            in1 => \N__31133\,
            in2 => \N__31121\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31112\,
            in2 => \N__31082\,
            in3 => \N__31100\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31073\,
            in2 => \N__31043\,
            in3 => \N__31061\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31031\,
            in2 => \N__31004\,
            in3 => \N__31019\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32609\,
            in2 => \N__30980\,
            in3 => \N__30995\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30971\,
            in2 => \N__30941\,
            in3 => \N__30956\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31364\,
            in2 => \N__31394\,
            in3 => \N__31379\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31358\,
            in1 => \N__31343\,
            in2 => \N__31331\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31319\,
            in1 => \N__32822\,
            in2 => \N__31304\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31295\,
            in1 => \N__31280\,
            in2 => \N__31271\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32597\,
            in2 => \N__32525\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31262\,
            in2 => \N__31250\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31232\,
            in2 => \N__31223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31208\,
            in2 => \N__31199\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31622\,
            in2 => \N__31613\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31601\,
            in2 => \N__31592\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31574\,
            in2 => \N__31562\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31547\,
            in2 => \N__31535\,
            in3 => \N__31499\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31496\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31489\,
            in2 => \_gnd_net_\,
            in3 => \N__35233\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31465\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35238\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35236\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31414\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__32503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35237\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32479\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__32455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35232\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35235\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32428\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010111"
        )
    port map (
            in0 => \N__32408\,
            in1 => \N__32384\,
            in2 => \N__32225\,
            in3 => \N__32031\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49038\,
            ce => 'H',
            sr => \N__48609\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33481\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49038\,
            ce => 'H',
            sr => \N__48609\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49038\,
            ce => 'H',
            sr => \N__48609\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31658\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32741\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32730\,
            in1 => \N__32708\,
            in2 => \_gnd_net_\,
            in3 => \N__34586\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49106\,
            ce => \N__34184\,
            sr => \N__48525\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34625\,
            in1 => \N__32662\,
            in2 => \_gnd_net_\,
            in3 => \N__32638\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34624\,
            in1 => \N__34767\,
            in2 => \_gnd_net_\,
            in3 => \N__34743\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32883\,
            in1 => \_gnd_net_\,
            in2 => \N__32930\,
            in3 => \N__34683\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49089\,
            ce => \N__34185\,
            sr => \N__48534\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34681\,
            in1 => \N__32769\,
            in2 => \_gnd_net_\,
            in3 => \N__32809\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49089\,
            ce => \N__34185\,
            sr => \N__48534\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32658\,
            in1 => \N__32642\,
            in2 => \_gnd_net_\,
            in3 => \N__34682\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49089\,
            ce => \N__34185\,
            sr => \N__48534\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__32562\,
            in1 => \N__32537\,
            in2 => \N__32585\,
            in3 => \N__32548\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__32580\,
            in1 => \N__32563\,
            in2 => \N__32549\,
            in3 => \N__32536\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34612\,
            in1 => \N__32887\,
            in2 => \_gnd_net_\,
            in3 => \N__32929\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32848\,
            in1 => \N__34613\,
            in2 => \_gnd_net_\,
            in3 => \N__32866\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34611\,
            in2 => \N__32852\,
            in3 => \N__32849\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49080\,
            ce => \N__34258\,
            sr => \N__48541\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32810\,
            in1 => \N__34610\,
            in2 => \_gnd_net_\,
            in3 => \N__32773\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33731\,
            in2 => \N__33692\,
            in3 => \N__33690\,
            lcout => \current_shift_inst.control_input_18\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33803\,
            in2 => \_gnd_net_\,
            in3 => \N__32753\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33797\,
            in2 => \_gnd_net_\,
            in3 => \N__32750\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33791\,
            in2 => \_gnd_net_\,
            in3 => \N__32747\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33785\,
            in2 => \_gnd_net_\,
            in3 => \N__32744\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33779\,
            in2 => \_gnd_net_\,
            in3 => \N__32957\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33773\,
            in2 => \_gnd_net_\,
            in3 => \N__32954\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33767\,
            in2 => \_gnd_net_\,
            in3 => \N__32951\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33761\,
            in2 => \_gnd_net_\,
            in3 => \N__32948\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33755\,
            in2 => \_gnd_net_\,
            in3 => \N__32945\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33122\,
            in2 => \_gnd_net_\,
            in3 => \N__32942\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36161\,
            in2 => \_gnd_net_\,
            in3 => \N__32939\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33671\,
            in2 => \_gnd_net_\,
            in3 => \N__32936\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44471\,
            in2 => \_gnd_net_\,
            in3 => \N__32933\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36098\,
            in1 => \N__36191\,
            in2 => \_gnd_net_\,
            in3 => \N__44470\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33107\,
            in2 => \_gnd_net_\,
            in3 => \N__33116\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33101\,
            in2 => \_gnd_net_\,
            in3 => \N__33071\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33068\,
            in3 => \N__33035\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33032\,
            in2 => \_gnd_net_\,
            in3 => \N__33023\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33020\,
            in2 => \_gnd_net_\,
            in3 => \N__32984\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32981\,
            in2 => \_gnd_net_\,
            in3 => \N__32972\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32969\,
            in2 => \_gnd_net_\,
            in3 => \N__32960\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33257\,
            in2 => \_gnd_net_\,
            in3 => \N__33248\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__49060\,
            ce => 'H',
            sr => \N__48565\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33245\,
            in2 => \_gnd_net_\,
            in3 => \N__33236\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33233\,
            in2 => \_gnd_net_\,
            in3 => \N__33224\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33221\,
            in2 => \_gnd_net_\,
            in3 => \N__33212\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33209\,
            in2 => \_gnd_net_\,
            in3 => \N__33200\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33197\,
            in2 => \_gnd_net_\,
            in3 => \N__33164\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33971\,
            in2 => \_gnd_net_\,
            in3 => \N__33161\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33986\,
            in2 => \_gnd_net_\,
            in3 => \N__33158\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33151\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49052\,
            ce => 'H',
            sr => \N__48574\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33507\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33465\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33432\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33405\,
            in2 => \_gnd_net_\,
            in3 => \N__35177\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33372\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__33342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35174\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33318\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33282\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__35881\,
            in1 => \N__34903\,
            in2 => \N__34888\,
            in3 => \N__33565\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49037\,
            ce => 'H',
            sr => \N__48590\
        );

    \phase_controller_inst2.state_ns_i_a2_1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35058\,
            in2 => \_gnd_net_\,
            in3 => \N__34818\,
            lcout => state_ns_i_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34902\,
            in2 => \_gnd_net_\,
            in3 => \N__33564\,
            lcout => \phase_controller_inst1.N_55\,
            ltout => \phase_controller_inst1.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__36336\,
            in1 => \N__39219\,
            in2 => \N__33662\,
            in3 => \N__33652\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49037\,
            ce => 'H',
            sr => \N__48590\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35239\,
            in2 => \_gnd_net_\,
            in3 => \N__33636\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__36337\,
            in1 => \N__39195\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__34796\,
            in1 => \N__34884\,
            in2 => \_gnd_net_\,
            in3 => \N__35872\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49026\,
            ce => 'H',
            sr => \N__48610\
        );

    \phase_controller_inst2.start_timer_hc_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__34837\,
            in1 => \N__33617\,
            in2 => \N__35804\,
            in3 => \N__33602\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49026\,
            ce => 'H',
            sr => \N__48610\
        );

    \phase_controller_inst1.T23_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__33583\,
            in1 => \N__35873\,
            in2 => \_gnd_net_\,
            in3 => \N__33571\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49021\,
            ce => 'H',
            sr => \N__48618\
        );

    \phase_controller_inst1.T45_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__33572\,
            in1 => \N__33535\,
            in2 => \_gnd_net_\,
            in3 => \N__39214\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49021\,
            ce => 'H',
            sr => \N__48618\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41023\,
            in1 => \N__40986\,
            in2 => \_gnd_net_\,
            in3 => \N__49336\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37049\,
            in2 => \_gnd_net_\,
            in3 => \N__35811\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35813\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49008\,
            ce => 'H',
            sr => \N__48656\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34975\,
            in2 => \_gnd_net_\,
            in3 => \N__35092\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__42165\,
            in1 => \N__44305\,
            in2 => \N__41411\,
            in3 => \N__44728\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44733\,
            in1 => \N__46646\,
            in2 => \N__41705\,
            in3 => \N__42163\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42161\,
            in1 => \N__44735\,
            in2 => \N__46328\,
            in3 => \N__39110\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44729\,
            in1 => \N__42166\,
            in2 => \N__44234\,
            in3 => \N__41542\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45694\,
            in1 => \N__44730\,
            in2 => \N__42319\,
            in3 => \N__41332\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44732\,
            in1 => \N__42162\,
            in2 => \N__46724\,
            in3 => \N__38980\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__42164\,
            in1 => \N__44731\,
            in2 => \N__41582\,
            in3 => \N__45170\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44734\,
            in1 => \N__46574\,
            in2 => \N__42320\,
            in3 => \N__38948\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33965\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49100\,
            ce => 'H',
            sr => \N__48529\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45479\,
            in1 => \N__41864\,
            in2 => \_gnd_net_\,
            in3 => \N__38911\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45478\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__35912\,
            in1 => \N__36152\,
            in2 => \_gnd_net_\,
            in3 => \N__44426\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33725\,
            in3 => \N__33691\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49092\,
            ce => 'H',
            sr => \N__48535\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44427\,
            lcout => \current_shift_inst.N_1326_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44429\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__44428\,
            in1 => \N__36143\,
            in2 => \_gnd_net_\,
            in3 => \N__35897\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__36134\,
            in1 => \N__36050\,
            in2 => \_gnd_net_\,
            in3 => \N__44462\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__44463\,
            in1 => \N__36125\,
            in2 => \_gnd_net_\,
            in3 => \N__36035\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36011\,
            in1 => \N__36116\,
            in2 => \_gnd_net_\,
            in3 => \N__44464\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__44465\,
            in1 => \N__35990\,
            in2 => \_gnd_net_\,
            in3 => \N__36236\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__35966\,
            in1 => \N__36227\,
            in2 => \_gnd_net_\,
            in3 => \N__44466\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__44467\,
            in1 => \N__35954\,
            in2 => \_gnd_net_\,
            in3 => \N__36218\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__35942\,
            in1 => \N__36209\,
            in2 => \_gnd_net_\,
            in3 => \N__44468\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__44469\,
            in1 => \N__35924\,
            in2 => \_gnd_net_\,
            in3 => \N__36200\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34772\,
            in1 => \N__34745\,
            in2 => \_gnd_net_\,
            in3 => \N__34687\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49073\,
            ce => \N__34155\,
            sr => \N__48546\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49452\,
            in1 => \N__35768\,
            in2 => \_gnd_net_\,
            in3 => \N__40214\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49066\,
            ce => \N__49982\,
            sr => \N__48554\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36300\,
            in1 => \N__39932\,
            in2 => \_gnd_net_\,
            in3 => \N__49453\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49066\,
            ce => \N__49982\,
            sr => \N__48554\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33982\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33951\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33912\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33867\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35651\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33825\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__35121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35217\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__34820\,
            in1 => \N__35105\,
            in2 => \N__34850\,
            in3 => \N__35088\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49053\,
            ce => 'H',
            sr => \N__48575\
        );

    \phase_controller_inst1.state_4_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35037\,
            in2 => \_gnd_net_\,
            in3 => \N__34819\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49053\,
            ce => 'H',
            sr => \N__48575\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__35002\,
            in1 => \N__34904\,
            in2 => \N__34982\,
            in3 => \N__34942\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49053\,
            ce => 'H',
            sr => \N__48575\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__35880\,
            in1 => \N__39167\,
            in2 => \N__34889\,
            in3 => \N__39253\,
            lcout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39279\,
            in1 => \N__40279\,
            in2 => \_gnd_net_\,
            in3 => \N__49429\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39166\,
            in2 => \_gnd_net_\,
            in3 => \N__39252\,
            lcout => \phase_controller_inst1.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__34836\,
            in1 => \N__34792\,
            in2 => \N__34781\,
            in3 => \N__50132\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49039\,
            ce => 'H',
            sr => \N__48591\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50133\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49039\,
            ce => 'H',
            sr => \N__48591\
        );

    \phase_controller_inst1.T12_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__35494\,
            in1 => \N__35871\,
            in2 => \_gnd_net_\,
            in3 => \N__39172\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49039\,
            ce => 'H',
            sr => \N__48591\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36259\,
            in1 => \N__40075\,
            in2 => \_gnd_net_\,
            in3 => \N__49546\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35573\,
            in1 => \N__40144\,
            in2 => \_gnd_net_\,
            in3 => \N__49547\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49031\,
            ce => \N__50031\,
            sr => \N__48601\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40211\,
            in2 => \_gnd_net_\,
            in3 => \N__40278\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__47095\,
            in1 => \N__49709\,
            in2 => \N__35483\,
            in3 => \N__35480\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43874\,
            in1 => \N__49418\,
            in2 => \_gnd_net_\,
            in3 => \N__40908\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__35650\,
            in1 => \N__35702\,
            in2 => \_gnd_net_\,
            in3 => \N__35680\,
            lcout => \current_shift_inst.timer_s1.N_168_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40001\,
            in1 => \N__40074\,
            in2 => \N__39920\,
            in3 => \N__40139\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35472\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__35540\,
            in1 => \N__35549\,
            in2 => \N__36491\,
            in3 => \N__36468\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__35548\,
            in1 => \N__36489\,
            in2 => \N__36470\,
            in3 => \N__35539\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49419\,
            in1 => \N__43499\,
            in2 => \_gnd_net_\,
            in3 => \N__39830\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49022\,
            ce => \N__48719\,
            sr => \N__48619\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43529\,
            in1 => \N__39860\,
            in2 => \_gnd_net_\,
            in3 => \N__49421\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49022\,
            ce => \N__48719\,
            sr => \N__48619\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40070\,
            in1 => \N__36260\,
            in2 => \_gnd_net_\,
            in3 => \N__49420\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49022\,
            ce => \N__48719\,
            sr => \N__48619\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__36405\,
            in1 => \N__36510\,
            in2 => \N__35522\,
            in3 => \N__35531\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__35530\,
            in1 => \N__36406\,
            in2 => \N__36512\,
            in3 => \N__35518\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48112\,
            in1 => \N__47595\,
            in2 => \_gnd_net_\,
            in3 => \N__49353\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49018\,
            ce => \N__48717\,
            sr => \N__48626\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47703\,
            in1 => \N__49350\,
            in2 => \_gnd_net_\,
            in3 => \N__47686\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49018\,
            ce => \N__48717\,
            sr => \N__48626\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49320\,
            in1 => \N__35568\,
            in2 => \_gnd_net_\,
            in3 => \N__40140\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47599\,
            in1 => \N__48107\,
            in2 => \_gnd_net_\,
            in3 => \N__49318\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__38309\,
            in1 => \N__35594\,
            in2 => \N__48023\,
            in3 => \N__41016\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__47707\,
            in1 => \_gnd_net_\,
            in2 => \N__35585\,
            in3 => \N__47679\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50197\,
            in1 => \N__50172\,
            in2 => \_gnd_net_\,
            in3 => \N__49321\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49319\,
            in1 => \N__35763\,
            in2 => \_gnd_net_\,
            in3 => \N__40212\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43840\,
            in1 => \N__49335\,
            in2 => \_gnd_net_\,
            in3 => \N__47809\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35646\,
            in2 => \_gnd_net_\,
            in3 => \N__35679\,
            lcout => \current_shift_inst.timer_s1.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36280\,
            in1 => \N__40002\,
            in2 => \_gnd_net_\,
            in3 => \N__49334\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49573\,
            in1 => \N__35569\,
            in2 => \_gnd_net_\,
            in3 => \N__40145\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49012\,
            ce => \N__48712\,
            sr => \N__48642\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__39280\,
            in1 => \_gnd_net_\,
            in2 => \N__49578\,
            in3 => \N__40280\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49012\,
            ce => \N__48712\,
            sr => \N__48642\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__35764\,
            in1 => \_gnd_net_\,
            in2 => \N__49579\,
            in3 => \N__40213\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49012\,
            ce => \N__48712\,
            sr => \N__48642\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49572\,
            in1 => \N__43836\,
            in2 => \_gnd_net_\,
            in3 => \N__47810\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49012\,
            ce => \N__48712\,
            sr => \N__48642\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49469\,
            in1 => \N__36276\,
            in2 => \_gnd_net_\,
            in3 => \N__40003\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49012\,
            ce => \N__48712\,
            sr => \N__48642\
        );

    \current_shift_inst.stop_timer_s1_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__35608\,
            in1 => \N__39229\,
            in2 => \N__35681\,
            in3 => \N__35700\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49011\,
            ce => 'H',
            sr => \N__48647\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000001100"
        )
    port map (
            in0 => \N__37067\,
            in1 => \N__35724\,
            in2 => \N__37277\,
            in3 => \N__37051\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49011\,
            ce => 'H',
            sr => \N__48647\
        );

    \current_shift_inst.start_timer_s1_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__35699\,
            in2 => \_gnd_net_\,
            in3 => \N__39228\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49011\,
            ce => 'H',
            sr => \N__48647\
        );

    \current_shift_inst.timer_s1.running_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__35701\,
            in1 => \N__35675\,
            in2 => \_gnd_net_\,
            in3 => \N__35645\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49011\,
            ce => 'H',
            sr => \N__48647\
        );

    \phase_controller_inst1.S1_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39230\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49011\,
            ce => 'H',
            sr => \N__48647\
        );

    \phase_controller_inst2.stoper_hc.running_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__37050\,
            in1 => \N__37066\,
            in2 => \N__35828\,
            in3 => \N__37273\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49009\,
            ce => 'H',
            sr => \N__48650\
        );

    \phase_controller_inst1.S2_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35885\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49009\,
            ce => 'H',
            sr => \N__48650\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__37048\,
            in1 => \N__35824\,
            in2 => \_gnd_net_\,
            in3 => \N__35812\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__38553\,
            in1 => \N__40889\,
            in2 => \N__38600\,
            in3 => \N__40959\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39594\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35777\,
            ce => 'H',
            sr => \N__48517\
        );

    \delay_measurement_inst.start_timer_hc_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39593\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35777\,
            ce => 'H',
            sr => \N__48517\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37622\,
            in2 => \N__37640\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37590\,
            in2 => \N__37205\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42213\,
            in2 => \N__37496\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37523\,
            in2 => \N__42387\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42217\,
            in2 => \N__37217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37544\,
            in2 => \N__42388\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42221\,
            in2 => \N__37178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37550\,
            in2 => \N__42389\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42225\,
            in2 => \N__37187\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37166\,
            in2 => \N__42390\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42229\,
            in2 => \N__37532\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38771\,
            in2 => \N__42391\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42233\,
            in2 => \N__38762\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38483\,
            in2 => \N__42392\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42237\,
            in2 => \N__37196\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38492\,
            in2 => \N__42393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42241\,
            in2 => \N__38726\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42245\,
            in2 => \N__37706\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42242\,
            in2 => \N__38714\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42246\,
            in2 => \N__39047\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42243\,
            in2 => \N__38750\,
            in3 => \N__35900\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42247\,
            in2 => \N__41894\,
            in3 => \N__35888\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42244\,
            in2 => \N__38738\,
            in3 => \N__36038\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42248\,
            in2 => \N__38699\,
            in3 => \N__36023\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42131\,
            in2 => \N__36020\,
            in3 => \N__35999\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35996\,
            in2 => \N__42303\,
            in3 => \N__35978\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42135\,
            in2 => \N__35975\,
            in3 => \N__35957\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37517\,
            in2 => \N__42304\,
            in3 => \N__35945\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42139\,
            in2 => \N__42530\,
            in3 => \N__35933\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35930\,
            in2 => \N__42305\,
            in3 => \N__35915\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42143\,
            in2 => \N__37724\,
            in3 => \N__36086\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__42144\,
            in1 => \N__44752\,
            in2 => \_gnd_net_\,
            in3 => \N__36083\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37615\,
            in2 => \N__37484\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43798\,
            in1 => \N__37583\,
            in2 => \N__37559\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42103\,
            in2 => \N__37508\,
            in3 => \N__43799\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36080\,
            in2 => \N__42296\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42107\,
            in2 => \N__36068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38504\,
            in2 => \N__42297\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42111\,
            in2 => \N__36059\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40844\,
            in2 => \N__42298\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42115\,
            in2 => \N__37685\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37781\,
            in2 => \N__42299\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42119\,
            in2 => \N__37793\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37775\,
            in2 => \N__42300\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42123\,
            in2 => \N__37715\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36107\,
            in2 => \N__42301\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42127\,
            in2 => \N__37694\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37730\,
            in2 => \N__42302\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42249\,
            in2 => \N__37811\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37754\,
            in2 => \N__42394\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42253\,
            in2 => \N__37748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37769\,
            in2 => \N__42395\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42257\,
            in2 => \N__37739\,
            in3 => \N__36146\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42485\,
            in2 => \N__42396\,
            in3 => \N__36137\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42261\,
            in2 => \N__37763\,
            in3 => \N__36128\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39056\,
            in2 => \N__42397\,
            in3 => \N__36119\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42306\,
            in2 => \N__37850\,
            in3 => \N__36110\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37835\,
            in2 => \N__42422\,
            in3 => \N__36230\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42310\,
            in2 => \N__37829\,
            in3 => \N__36221\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37802\,
            in2 => \N__42423\,
            in3 => \N__36212\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42314\,
            in2 => \N__37862\,
            in3 => \N__36203\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37841\,
            in2 => \N__42424\,
            in3 => \N__36194\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42318\,
            in2 => \N__37820\,
            in3 => \N__36182\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__42497\,
            in1 => \N__44461\,
            in2 => \N__36179\,
            in3 => \N__36164\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36304\,
            in1 => \N__39928\,
            in2 => \_gnd_net_\,
            in3 => \N__49580\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48680\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__39215\,
            in1 => \N__39168\,
            in2 => \N__36341\,
            in3 => \N__39254\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49054\,
            ce => 'H',
            sr => \N__48576\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49479\,
            in1 => \N__47378\,
            in2 => \_gnd_net_\,
            in3 => \N__47396\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49047\,
            ce => \N__48722\,
            sr => \N__48584\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36308\,
            in1 => \N__39927\,
            in2 => \_gnd_net_\,
            in3 => \N__49481\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49047\,
            ce => \N__48722\,
            sr => \N__48584\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47850\,
            in1 => \N__49480\,
            in2 => \_gnd_net_\,
            in3 => \N__46913\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49047\,
            ce => \N__48722\,
            sr => \N__48584\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36284\,
            in1 => \N__40004\,
            in2 => \_gnd_net_\,
            in3 => \N__49550\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49040\,
            ce => \N__50027\,
            sr => \N__48592\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49548\,
            in1 => \N__41027\,
            in2 => \_gnd_net_\,
            in3 => \N__40990\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49040\,
            ce => \N__50027\,
            sr => \N__48592\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36255\,
            in1 => \N__40076\,
            in2 => \_gnd_net_\,
            in3 => \N__49549\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49040\,
            ce => \N__50027\,
            sr => \N__48592\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37247\,
            in2 => \N__37466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37417\,
            in1 => \N__36538\,
            in2 => \_gnd_net_\,
            in3 => \N__36239\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__37425\,
            in1 => \N__36805\,
            in2 => \N__37454\,
            in3 => \N__36389\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37418\,
            in1 => \N__36781\,
            in2 => \_gnd_net_\,
            in3 => \N__36386\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37426\,
            in1 => \N__36754\,
            in2 => \_gnd_net_\,
            in3 => \N__36383\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37419\,
            in1 => \N__36730\,
            in2 => \_gnd_net_\,
            in3 => \N__36380\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37427\,
            in1 => \N__36700\,
            in2 => \_gnd_net_\,
            in3 => \N__36377\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37420\,
            in1 => \N__36670\,
            in2 => \_gnd_net_\,
            in3 => \N__36374\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49032\,
            ce => 'H',
            sr => \N__48602\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37431\,
            in1 => \N__36640\,
            in2 => \_gnd_net_\,
            in3 => \N__36371\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37413\,
            in1 => \N__37003\,
            in2 => \_gnd_net_\,
            in3 => \N__36368\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37428\,
            in1 => \N__36961\,
            in2 => \_gnd_net_\,
            in3 => \N__36365\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37414\,
            in1 => \N__36925\,
            in2 => \_gnd_net_\,
            in3 => \N__36431\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37429\,
            in1 => \N__36892\,
            in2 => \_gnd_net_\,
            in3 => \N__36428\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37415\,
            in1 => \N__36856\,
            in2 => \_gnd_net_\,
            in3 => \N__36425\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37430\,
            in1 => \N__36829\,
            in2 => \_gnd_net_\,
            in3 => \N__36422\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37416\,
            in1 => \N__38261\,
            in2 => \_gnd_net_\,
            in3 => \N__36419\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49027\,
            ce => 'H',
            sr => \N__48611\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37421\,
            in1 => \N__38241\,
            in2 => \_gnd_net_\,
            in3 => \N__36416\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37432\,
            in1 => \N__38665\,
            in2 => \_gnd_net_\,
            in3 => \N__36413\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37422\,
            in1 => \N__38641\,
            in2 => \_gnd_net_\,
            in3 => \N__36410\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37433\,
            in1 => \N__36407\,
            in2 => \_gnd_net_\,
            in3 => \N__36392\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37423\,
            in1 => \N__36511\,
            in2 => \_gnd_net_\,
            in3 => \N__36494\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37434\,
            in1 => \N__36490\,
            in2 => \_gnd_net_\,
            in3 => \N__36473\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37424\,
            in1 => \N__36469\,
            in2 => \_gnd_net_\,
            in3 => \N__36452\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37435\,
            in1 => \N__36579\,
            in2 => \_gnd_net_\,
            in3 => \N__36449\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49023\,
            ce => 'H',
            sr => \N__48620\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37402\,
            in1 => \N__36599\,
            in2 => \_gnd_net_\,
            in3 => \N__36446\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37406\,
            in1 => \N__38474\,
            in2 => \_gnd_net_\,
            in3 => \N__36443\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37403\,
            in1 => \N__38451\,
            in2 => \_gnd_net_\,
            in3 => \N__36440\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37407\,
            in1 => \N__38405\,
            in2 => \_gnd_net_\,
            in3 => \N__36437\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37404\,
            in1 => \N__38389\,
            in2 => \_gnd_net_\,
            in3 => \N__36434\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37408\,
            in1 => \N__38543\,
            in2 => \_gnd_net_\,
            in3 => \N__36617\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37405\,
            in1 => \N__38582\,
            in2 => \_gnd_net_\,
            in3 => \N__36614\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49019\,
            ce => 'H',
            sr => \N__48627\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__36598\,
            in1 => \N__36580\,
            in2 => \N__36563\,
            in3 => \N__36611\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36610\,
            in1 => \N__36597\,
            in2 => \N__36584\,
            in3 => \N__36559\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47918\,
            in1 => \N__47959\,
            in2 => \_gnd_net_\,
            in3 => \N__49352\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49014\,
            ce => \N__48714\,
            sr => \N__48633\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49351\,
            in1 => \N__50193\,
            in2 => \_gnd_net_\,
            in3 => \N__50177\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49014\,
            ce => \N__48714\,
            sr => \N__48633\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__38299\,
            in1 => \N__38473\,
            in2 => \N__38455\,
            in3 => \N__38341\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38324\,
            in2 => \N__36551\,
            in3 => \N__37243\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36542\,
            in1 => \N__38612\,
            in2 => \N__36524\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36791\,
            in2 => \N__38351\,
            in3 => \N__36809\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38330\,
            in2 => \N__36767\,
            in3 => \N__36785\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49157\,
            in2 => \N__36740\,
            in3 => \N__36758\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38357\,
            in2 => \N__36716\,
            in3 => \N__36731\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36707\,
            in2 => \N__36686\,
            in3 => \N__36701\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36677\,
            in2 => \N__36656\,
            in3 => \N__36671\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36647\,
            in2 => \N__36626\,
            in3 => \N__36641\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37004\,
            in1 => \N__36989\,
            in2 => \N__36977\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36968\,
            in2 => \N__36947\,
            in3 => \N__36962\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36911\,
            in2 => \N__36938\,
            in3 => \N__36926\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36878\,
            in2 => \N__36905\,
            in3 => \N__36896\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36872\,
            in2 => \N__36842\,
            in3 => \N__36857\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36830\,
            in1 => \N__36815\,
            in2 => \N__40856\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38273\,
            in2 => \N__38225\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38618\,
            in2 => \N__38684\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37160\,
            in2 => \N__37148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37133\,
            in2 => \N__37121\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37103\,
            in2 => \N__37094\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37082\,
            in2 => \N__38429\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38414\,
            in2 => \N__38372\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38606\,
            in2 => \N__38519\,
            in3 => \N__37073\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37070\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__38515\,
            in1 => \N__37055\,
            in2 => \N__37019\,
            in3 => \N__37010\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37469\,
            in3 => \N__37268\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37267\,
            in2 => \_gnd_net_\,
            in3 => \N__37285\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__37409\,
            in1 => \N__37286\,
            in2 => \N__37242\,
            in3 => \N__37269\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49010\,
            ce => 'H',
            sr => \N__48651\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44678\,
            in1 => \N__42452\,
            in2 => \N__41543\,
            in3 => \N__44230\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41384\,
            in1 => \N__44677\,
            in2 => \N__37598\,
            in3 => \N__41362\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__42438\,
            in1 => \N__44598\,
            in2 => \N__41207\,
            in3 => \N__46252\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44595\,
            in1 => \N__42443\,
            in2 => \N__45562\,
            in3 => \N__41308\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__42441\,
            in1 => \N__41333\,
            in2 => \N__45698\,
            in3 => \N__44593\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44596\,
            in1 => \N__42444\,
            in2 => \N__38912\,
            in3 => \N__45477\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__42442\,
            in1 => \N__44594\,
            in2 => \N__41432\,
            in3 => \N__45626\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44592\,
            in1 => \N__42440\,
            in2 => \N__44155\,
            in3 => \N__41515\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42437\,
            in1 => \N__44597\,
            in2 => \N__45404\,
            in3 => \N__41753\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44591\,
            in1 => \N__42439\,
            in2 => \N__44309\,
            in3 => \N__41407\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42325\,
            in1 => \N__44556\,
            in2 => \N__46505\,
            in3 => \N__41606\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47135\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49130\,
            ce => \N__47168\,
            sr => \N__48518\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42326\,
            in1 => \N__44552\,
            in2 => \N__44366\,
            in3 => \N__41182\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__41183\,
            in1 => \N__44362\,
            in2 => \N__44657\,
            in3 => \N__42327\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37667\,
            in1 => \N__44551\,
            in2 => \_gnd_net_\,
            in3 => \N__37676\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38826\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37666\,
            in2 => \N__37670\,
            in3 => \N__44550\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44393\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49123\,
            ce => \N__47166\,
            sr => \N__48519\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37664\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__37665\,
            in1 => \_gnd_net_\,
            in2 => \N__37646\,
            in3 => \N__41847\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__44890\,
            in1 => \N__43765\,
            in2 => \_gnd_net_\,
            in3 => \N__37604\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44891\,
            in2 => \N__37643\,
            in3 => \N__37636\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47134\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49123\,
            ce => \N__47166\,
            sr => \N__48519\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41848\,
            in1 => \N__45312\,
            in2 => \_gnd_net_\,
            in3 => \N__38871\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44658\,
            in1 => \N__41380\,
            in2 => \N__37591\,
            in3 => \N__41352\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49116\,
            ce => \N__47163\,
            sr => \N__48522\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41351\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44659\,
            in2 => \_gnd_net_\,
            in3 => \N__39075\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__44660\,
            in1 => \N__42160\,
            in2 => \N__39080\,
            in3 => \N__43800\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42182\,
            in1 => \N__44665\,
            in2 => \N__45247\,
            in3 => \N__41491\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44667\,
            in1 => \N__46037\,
            in2 => \N__42323\,
            in3 => \N__41677\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42183\,
            in1 => \N__44666\,
            in2 => \N__46256\,
            in3 => \N__41203\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44668\,
            in1 => \N__46320\,
            in2 => \_gnd_net_\,
            in3 => \N__39102\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42184\,
            in1 => \N__44661\,
            in2 => \N__45563\,
            in3 => \N__41309\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44663\,
            in1 => \N__45403\,
            in2 => \N__42321\,
            in3 => \N__41749\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45476\,
            in1 => \N__44662\,
            in2 => \N__42324\,
            in3 => \N__38904\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44664\,
            in1 => \N__45322\,
            in2 => \N__42322\,
            in3 => \N__38872\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44713\,
            in1 => \N__45895\,
            in2 => \N__42469\,
            in3 => \N__42548\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__41468\,
            in1 => \N__42407\,
            in2 => \N__46865\,
            in3 => \N__44715\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44711\,
            in1 => \N__46036\,
            in2 => \N__42468\,
            in3 => \N__41678\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__45967\,
            in1 => \N__44712\,
            in2 => \N__41660\,
            in3 => \N__42416\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44714\,
            in1 => \N__45823\,
            in2 => \N__42467\,
            in3 => \N__41728\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__41168\,
            in1 => \N__44710\,
            in2 => \N__46193\,
            in3 => \N__42412\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44717\,
            in1 => \N__46409\,
            in2 => \N__42466\,
            in3 => \N__42514\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__46720\,
            in1 => \N__44716\,
            in2 => \N__38987\,
            in3 => \N__42411\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__39106\,
            in1 => \N__46324\,
            in2 => \N__42471\,
            in3 => \N__44723\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44720\,
            in1 => \N__46645\,
            in2 => \N__42472\,
            in3 => \N__41698\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__42431\,
            in1 => \N__38941\,
            in2 => \N__46570\,
            in3 => \N__44721\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__44724\,
            in1 => \N__42433\,
            in2 => \N__39079\,
            in3 => \N__43807\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46563\,
            in1 => \N__44719\,
            in2 => \_gnd_net_\,
            in3 => \N__38940\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44718\,
            in1 => \N__42432\,
            in2 => \N__46111\,
            in3 => \N__42575\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__41602\,
            in1 => \N__46501\,
            in2 => \N__42470\,
            in3 => \N__44722\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38125\,
            in1 => \N__44385\,
            in2 => \_gnd_net_\,
            in3 => \N__37796\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38117\,
            in1 => \N__44328\,
            in2 => \_gnd_net_\,
            in3 => \N__37889\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_2_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38126\,
            in1 => \N__44248\,
            in2 => \_gnd_net_\,
            in3 => \N__37886\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38118\,
            in1 => \N__44170\,
            in2 => \_gnd_net_\,
            in3 => \N__37883\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_4_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38127\,
            in1 => \N__45714\,
            in2 => \_gnd_net_\,
            in3 => \N__37880\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_5_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38119\,
            in1 => \N__45640\,
            in2 => \_gnd_net_\,
            in3 => \N__37877\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_6_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38128\,
            in1 => \N__45577\,
            in2 => \_gnd_net_\,
            in3 => \N__37874\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_7_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38120\,
            in1 => \N__45493\,
            in2 => \_gnd_net_\,
            in3 => \N__37871\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__49083\,
            ce => \N__38002\,
            sr => \N__48542\
        );

    \current_shift_inst.timer_s1.counter_8_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38124\,
            in1 => \N__45426\,
            in2 => \_gnd_net_\,
            in3 => \N__37868\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_9_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38132\,
            in1 => \N__45345\,
            in2 => \_gnd_net_\,
            in3 => \N__37865\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_10_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38121\,
            in1 => \N__45264\,
            in2 => \_gnd_net_\,
            in3 => \N__37916\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_11_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38129\,
            in1 => \N__45186\,
            in2 => \_gnd_net_\,
            in3 => \N__37913\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_12_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38122\,
            in1 => \N__46272\,
            in2 => \_gnd_net_\,
            in3 => \N__37910\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_13_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38130\,
            in1 => \N__46207\,
            in2 => \_gnd_net_\,
            in3 => \N__37907\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_14_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38123\,
            in1 => \N__46128\,
            in2 => \_gnd_net_\,
            in3 => \N__37904\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_15_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38131\,
            in1 => \N__46051\,
            in2 => \_gnd_net_\,
            in3 => \N__37901\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__49074\,
            ce => \N__38003\,
            sr => \N__48547\
        );

    \current_shift_inst.timer_s1.counter_16_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38085\,
            in1 => \N__45987\,
            in2 => \_gnd_net_\,
            in3 => \N__37898\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_17_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38095\,
            in1 => \N__45912\,
            in2 => \_gnd_net_\,
            in3 => \N__37895\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_18_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38086\,
            in1 => \N__45843\,
            in2 => \_gnd_net_\,
            in3 => \N__37892\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_19_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38096\,
            in1 => \N__45771\,
            in2 => \_gnd_net_\,
            in3 => \N__37943\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_20_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38087\,
            in1 => \N__46879\,
            in2 => \_gnd_net_\,
            in3 => \N__37940\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_21_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38097\,
            in1 => \N__46810\,
            in2 => \_gnd_net_\,
            in3 => \N__37937\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_22_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38088\,
            in1 => \N__46738\,
            in2 => \_gnd_net_\,
            in3 => \N__37934\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_23_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38098\,
            in1 => \N__46660\,
            in2 => \_gnd_net_\,
            in3 => \N__37931\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__49067\,
            ce => \N__38001\,
            sr => \N__48555\
        );

    \current_shift_inst.timer_s1.counter_24_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38089\,
            in1 => \N__46590\,
            in2 => \_gnd_net_\,
            in3 => \N__37928\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__49061\,
            ce => \N__37991\,
            sr => \N__48566\
        );

    \current_shift_inst.timer_s1.counter_25_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38093\,
            in1 => \N__46521\,
            in2 => \_gnd_net_\,
            in3 => \N__37925\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__49061\,
            ce => \N__37991\,
            sr => \N__48566\
        );

    \current_shift_inst.timer_s1.counter_26_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38090\,
            in1 => \N__46431\,
            in2 => \_gnd_net_\,
            in3 => \N__37922\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__49061\,
            ce => \N__37991\,
            sr => \N__48566\
        );

    \current_shift_inst.timer_s1.counter_27_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38094\,
            in1 => \N__46344\,
            in2 => \_gnd_net_\,
            in3 => \N__37919\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__49061\,
            ce => \N__37991\,
            sr => \N__48566\
        );

    \current_shift_inst.timer_s1.counter_28_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38091\,
            in1 => \N__46450\,
            in2 => \_gnd_net_\,
            in3 => \N__38135\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__49061\,
            ce => \N__37991\,
            sr => \N__48566\
        );

    \current_shift_inst.timer_s1.counter_29_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__46369\,
            in1 => \N__38092\,
            in2 => \_gnd_net_\,
            in3 => \N__38006\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49061\,
            ce => \N__37991\,
            sr => \N__48566\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39517\,
            in1 => \N__39789\,
            in2 => \_gnd_net_\,
            in3 => \N__37964\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39521\,
            in1 => \N__39732\,
            in2 => \_gnd_net_\,
            in3 => \N__37961\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39518\,
            in1 => \N__40353\,
            in2 => \_gnd_net_\,
            in3 => \N__37958\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39522\,
            in1 => \N__40321\,
            in2 => \_gnd_net_\,
            in3 => \N__37955\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39519\,
            in1 => \N__40299\,
            in2 => \_gnd_net_\,
            in3 => \N__37952\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39523\,
            in1 => \N__40230\,
            in2 => \_gnd_net_\,
            in3 => \N__37949\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39520\,
            in1 => \N__40161\,
            in2 => \_gnd_net_\,
            in3 => \N__37946\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39524\,
            in1 => \N__40092\,
            in2 => \_gnd_net_\,
            in3 => \N__38162\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__49055\,
            ce => \N__39569\,
            sr => \N__48577\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39504\,
            in1 => \N__40023\,
            in2 => \_gnd_net_\,
            in3 => \N__38159\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39508\,
            in1 => \N__39951\,
            in2 => \_gnd_net_\,
            in3 => \N__38156\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39501\,
            in1 => \N__40596\,
            in2 => \_gnd_net_\,
            in3 => \N__38153\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39505\,
            in1 => \N__40575\,
            in2 => \_gnd_net_\,
            in3 => \N__38150\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39502\,
            in1 => \N__40551\,
            in2 => \_gnd_net_\,
            in3 => \N__38147\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39506\,
            in1 => \N__40524\,
            in2 => \_gnd_net_\,
            in3 => \N__38144\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39503\,
            in1 => \N__40494\,
            in2 => \_gnd_net_\,
            in3 => \N__38141\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39507\,
            in1 => \N__40467\,
            in2 => \_gnd_net_\,
            in3 => \N__38138\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__49048\,
            ce => \N__39574\,
            sr => \N__48585\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39509\,
            in1 => \N__40440\,
            in2 => \_gnd_net_\,
            in3 => \N__38189\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39536\,
            in1 => \N__40407\,
            in2 => \_gnd_net_\,
            in3 => \N__38186\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39510\,
            in1 => \N__40377\,
            in2 => \_gnd_net_\,
            in3 => \N__38183\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39537\,
            in1 => \N__40827\,
            in2 => \_gnd_net_\,
            in3 => \N__38180\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39511\,
            in1 => \N__40803\,
            in2 => \_gnd_net_\,
            in3 => \N__38177\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39538\,
            in1 => \N__40777\,
            in2 => \_gnd_net_\,
            in3 => \N__38174\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39512\,
            in1 => \N__40747\,
            in2 => \_gnd_net_\,
            in3 => \N__38171\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39539\,
            in1 => \N__40717\,
            in2 => \_gnd_net_\,
            in3 => \N__38168\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__49041\,
            ce => \N__39570\,
            sr => \N__48593\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39513\,
            in1 => \N__40692\,
            in2 => \_gnd_net_\,
            in3 => \N__38165\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__49033\,
            ce => \N__39575\,
            sr => \N__48603\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39534\,
            in1 => \N__40662\,
            in2 => \_gnd_net_\,
            in3 => \N__38288\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__49033\,
            ce => \N__39575\,
            sr => \N__48603\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39514\,
            in1 => \N__40620\,
            in2 => \_gnd_net_\,
            in3 => \N__38285\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__49033\,
            ce => \N__39575\,
            sr => \N__48603\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39535\,
            in1 => \N__41121\,
            in2 => \_gnd_net_\,
            in3 => \N__38282\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__49033\,
            ce => \N__39575\,
            sr => \N__48603\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39515\,
            in1 => \N__40639\,
            in2 => \_gnd_net_\,
            in3 => \N__38279\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__49033\,
            ce => \N__39575\,
            sr => \N__48603\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__41140\,
            in1 => \N__39516\,
            in2 => \_gnd_net_\,
            in3 => \N__38276\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49033\,
            ce => \N__39575\,
            sr => \N__48603\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__38259\,
            in1 => \N__38242\,
            in2 => \N__38201\,
            in3 => \N__38210\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__38209\,
            in1 => \N__38260\,
            in2 => \N__38246\,
            in3 => \N__38197\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49742\,
            in1 => \N__49769\,
            in2 => \_gnd_net_\,
            in3 => \N__49576\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49028\,
            ce => \N__48720\,
            sr => \N__48612\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49574\,
            in1 => \N__48172\,
            in2 => \_gnd_net_\,
            in3 => \N__47006\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49028\,
            ce => \N__48720\,
            sr => \N__48612\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49575\,
            in1 => \N__47250\,
            in2 => \_gnd_net_\,
            in3 => \N__47227\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49028\,
            ce => \N__48720\,
            sr => \N__48612\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39710\,
            in1 => \N__47756\,
            in2 => \N__39771\,
            in3 => \N__47225\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__50258\,
            in1 => \_gnd_net_\,
            in2 => \N__38312\,
            in3 => \N__43583\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49024\,
            ce => \N__41094\,
            sr => \N__48621\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49024\,
            ce => \N__41094\,
            sr => \N__48621\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47254\,
            in1 => \N__47226\,
            in2 => \_gnd_net_\,
            in3 => \N__49424\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47757\,
            in1 => \N__49425\,
            in2 => \_gnd_net_\,
            in3 => \N__47190\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39764\,
            in1 => \N__39330\,
            in2 => \_gnd_net_\,
            in3 => \N__49423\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49422\,
            in1 => \N__39303\,
            in2 => \_gnd_net_\,
            in3 => \N__39711\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__38300\,
            in1 => \N__38472\,
            in2 => \N__38456\,
            in3 => \N__38342\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__40864\,
            in1 => \N__40930\,
            in2 => \N__38390\,
            in3 => \N__38403\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__38404\,
            in1 => \N__40865\,
            in2 => \N__40931\,
            in3 => \N__38388\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43558\,
            in1 => \N__43584\,
            in2 => \_gnd_net_\,
            in3 => \N__49534\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47090\,
            in1 => \N__47041\,
            in2 => \_gnd_net_\,
            in3 => \N__49628\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49015\,
            ce => \N__48715\,
            sr => \N__48634\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47501\,
            in1 => \N__48149\,
            in2 => \_gnd_net_\,
            in3 => \N__49625\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49015\,
            ce => \N__48715\,
            sr => \N__48634\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49624\,
            in1 => \N__39334\,
            in2 => \_gnd_net_\,
            in3 => \N__39773\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49015\,
            ce => \N__48715\,
            sr => \N__48634\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50260\,
            in1 => \N__50236\,
            in2 => \_gnd_net_\,
            in3 => \N__49626\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49015\,
            ce => \N__48715\,
            sr => \N__48634\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39307\,
            in1 => \N__39716\,
            in2 => \_gnd_net_\,
            in3 => \N__49627\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49015\,
            ce => \N__48715\,
            sr => \N__48634\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100100010"
        )
    port map (
            in0 => \N__38627\,
            in1 => \N__38650\,
            in2 => \N__38675\,
            in3 => \N__41036\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__41035\,
            in1 => \N__38674\,
            in2 => \N__38651\,
            in3 => \N__38626\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47191\,
            in1 => \N__47764\,
            in2 => \_gnd_net_\,
            in3 => \N__49577\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49013\,
            ce => \N__48713\,
            sr => \N__48638\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101110001"
        )
    port map (
            in0 => \N__40961\,
            in1 => \N__38557\,
            in2 => \N__38599\,
            in3 => \N__40888\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__40887\,
            in1 => \N__38592\,
            in2 => \N__38558\,
            in3 => \N__40960\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__39396\,
            in1 => \N__39610\,
            in2 => \_gnd_net_\,
            in3 => \N__39379\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49140\,
            ce => 'H',
            sr => \N__48516\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44620\,
            in1 => \N__42451\,
            in2 => \N__44156\,
            in3 => \N__41516\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41167\,
            in1 => \N__44624\,
            in2 => \N__42473\,
            in3 => \N__46183\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44623\,
            in1 => \N__42447\,
            in2 => \N__45169\,
            in3 => \N__41572\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41863\,
            in1 => \N__46716\,
            in2 => \_gnd_net_\,
            in3 => \N__38973\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44621\,
            in1 => \N__42445\,
            in2 => \N__45323\,
            in3 => \N__38876\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42446\,
            in1 => \N__44622\,
            in2 => \N__45248\,
            in3 => \N__41495\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44222\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42459\,
            in1 => \N__44707\,
            in2 => \N__45827\,
            in3 => \N__41732\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45620\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41467\,
            in1 => \N__44708\,
            in2 => \N__42474\,
            in3 => \N__46861\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44705\,
            in1 => \N__42460\,
            in2 => \N__46112\,
            in3 => \N__42571\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42461\,
            in1 => \N__44706\,
            in2 => \N__45971\,
            in3 => \N__41653\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41627\,
            in1 => \N__44709\,
            in2 => \N__42475\,
            in3 => \N__46795\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38834\,
            in2 => \N__38827\,
            in3 => \N__38828\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41474\,
            in2 => \_gnd_net_\,
            in3 => \N__38804\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41444\,
            in2 => \_gnd_net_\,
            in3 => \N__38801\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38798\,
            in2 => \_gnd_net_\,
            in3 => \N__38792\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41711\,
            in2 => \_gnd_net_\,
            in3 => \N__38789\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41438\,
            in2 => \_gnd_net_\,
            in3 => \N__38786\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38783\,
            in2 => \_gnd_net_\,
            in3 => \N__38777\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41549\,
            in2 => \_gnd_net_\,
            in3 => \N__38774\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38924\,
            in2 => \_gnd_net_\,
            in3 => \N__38882\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42662\,
            in3 => \N__38879\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42632\,
            in3 => \N__38855\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42620\,
            in2 => \_gnd_net_\,
            in3 => \N__38852\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41633\,
            in2 => \_gnd_net_\,
            in3 => \N__38849\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42650\,
            in2 => \_gnd_net_\,
            in3 => \N__38846\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42596\,
            in2 => \_gnd_net_\,
            in3 => \N__38843\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39620\,
            in2 => \_gnd_net_\,
            in3 => \N__38840\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39023\,
            in2 => \_gnd_net_\,
            in3 => \N__38837\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42671\,
            in2 => \_gnd_net_\,
            in3 => \N__39005\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42641\,
            in2 => \_gnd_net_\,
            in3 => \N__39002\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42800\,
            in2 => \_gnd_net_\,
            in3 => \N__38999\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42791\,
            in3 => \N__38996\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42818\,
            in2 => \_gnd_net_\,
            in3 => \N__38993\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42608\,
            in3 => \N__38990\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42779\,
            in2 => \_gnd_net_\,
            in3 => \N__38954\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42767\,
            in2 => \_gnd_net_\,
            in3 => \N__38951\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39014\,
            in3 => \N__38927\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42809\,
            in2 => \_gnd_net_\,
            in3 => \N__39116\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39029\,
            in2 => \_gnd_net_\,
            in3 => \N__39113\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42584\,
            in2 => \_gnd_net_\,
            in3 => \N__39086\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39083\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__42420\,
            in1 => \N__44759\,
            in2 => \N__46796\,
            in3 => \N__41623\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44758\,
            in1 => \N__42421\,
            in2 => \N__45896\,
            in3 => \N__42547\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46406\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46028\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46562\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46094\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__39380\,
            in1 => \N__39407\,
            in2 => \_gnd_net_\,
            in3 => \N__39611\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39405\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39375\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39338\,
            in1 => \N__39772\,
            in2 => \_gnd_net_\,
            in3 => \N__49582\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49075\,
            ce => \N__49952\,
            sr => \N__48548\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39715\,
            in1 => \N__39308\,
            in2 => \_gnd_net_\,
            in3 => \N__49583\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49075\,
            ce => \N__49952\,
            sr => \N__48548\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49581\,
            in1 => \N__39281\,
            in2 => \_gnd_net_\,
            in3 => \N__40277\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49075\,
            ce => \N__49952\,
            sr => \N__48548\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001101000000"
        )
    port map (
            in0 => \N__43103\,
            in1 => \N__39670\,
            in2 => \N__50108\,
            in3 => \N__39251\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49068\,
            ce => 'H',
            sr => \N__48556\
        );

    \phase_controller_inst1.T01_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__39127\,
            in1 => \N__39227\,
            in2 => \_gnd_net_\,
            in3 => \N__39173\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49068\,
            ce => 'H',
            sr => \N__48556\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__39669\,
            in1 => \N__39878\,
            in2 => \N__43091\,
            in3 => \N__50052\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49068\,
            ce => 'H',
            sr => \N__48556\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__39679\,
            in1 => \N__50134\,
            in2 => \_gnd_net_\,
            in3 => \N__50098\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39683\,
            in3 => \N__39873\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__39680\,
            in1 => \N__43102\,
            in2 => \N__39671\,
            in3 => \N__50099\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49062\,
            ce => 'H',
            sr => \N__48567\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39665\,
            in2 => \_gnd_net_\,
            in3 => \N__39874\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__39635\,
            in1 => \N__39650\,
            in2 => \N__43703\,
            in3 => \N__43734\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__39649\,
            in1 => \N__39633\,
            in2 => \N__43735\,
            in3 => \N__43698\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__40915\,
            in1 => \N__43873\,
            in2 => \N__49623\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49056\,
            ce => \N__49994\,
            sr => \N__48578\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__39648\,
            in1 => \N__39634\,
            in2 => \N__43736\,
            in3 => \N__43699\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__50101\,
            in1 => \N__43126\,
            in2 => \N__39623\,
            in3 => \N__43115\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__39839\,
            in1 => \N__39809\,
            in2 => \N__43463\,
            in3 => \N__43440\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__39808\,
            in1 => \N__43461\,
            in2 => \N__43442\,
            in3 => \N__39838\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43524\,
            in1 => \N__39856\,
            in2 => \_gnd_net_\,
            in3 => \N__49530\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => \elapsed_time_ns_1_RNI14DN9_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49533\,
            in1 => \_gnd_net_\,
            in2 => \N__39842\,
            in3 => \N__43525\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49049\,
            ce => \N__50006\,
            sr => \N__48586\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43497\,
            in1 => \N__39823\,
            in2 => \_gnd_net_\,
            in3 => \N__49531\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49532\,
            in1 => \_gnd_net_\,
            in2 => \N__39812\,
            in3 => \N__43498\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49049\,
            ce => \N__50006\,
            sr => \N__48586\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40354\,
            in2 => \N__39800\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39739\,
            in2 => \N__40333\,
            in3 => \N__39686\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40355\,
            in2 => \N__40304\,
            in3 => \N__40337\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40231\,
            in2 => \N__40334\,
            in3 => \N__40307\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40303\,
            in2 => \N__40168\,
            in3 => \N__40235\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40232\,
            in2 => \N__40099\,
            in3 => \N__40172\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40024\,
            in2 => \N__40169\,
            in3 => \N__40103\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39952\,
            in2 => \N__40100\,
            in3 => \N__40034\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49042\,
            ce => \N__41087\,
            sr => \N__48594\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40597\,
            in2 => \N__40031\,
            in3 => \N__39962\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40576\,
            in2 => \N__39959\,
            in3 => \N__39881\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40598\,
            in2 => \N__40556\,
            in3 => \N__40580\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40577\,
            in2 => \N__40529\,
            in3 => \N__40559\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40555\,
            in2 => \N__40501\,
            in3 => \N__40532\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40528\,
            in2 => \N__40474\,
            in3 => \N__40505\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40441\,
            in2 => \N__40502\,
            in3 => \N__40478\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40414\,
            in2 => \N__40475\,
            in3 => \N__40451\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49034\,
            ce => \N__41083\,
            sr => \N__48604\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40378\,
            in2 => \N__40448\,
            in3 => \N__40421\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40828\,
            in2 => \N__40418\,
            in3 => \N__40385\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40804\,
            in2 => \N__40382\,
            in3 => \N__40358\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40783\,
            in2 => \N__40832\,
            in3 => \N__40808\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40805\,
            in2 => \N__40759\,
            in3 => \N__40787\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40784\,
            in2 => \N__40729\,
            in3 => \N__40763\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40693\,
            in2 => \N__40760\,
            in3 => \N__40733\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40663\,
            in2 => \N__40730\,
            in3 => \N__40703\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49029\,
            ce => \N__41095\,
            sr => \N__48613\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40621\,
            in2 => \N__40700\,
            in3 => \N__40673\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49025\,
            ce => \N__41096\,
            sr => \N__48622\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41122\,
            in2 => \N__40670\,
            in3 => \N__40643\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49025\,
            ce => \N__41096\,
            sr => \N__48622\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40640\,
            in2 => \N__40625\,
            in3 => \N__40601\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49025\,
            ce => \N__41096\,
            sr => \N__48622\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41144\,
            in2 => \N__41126\,
            in3 => \N__41102\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49025\,
            ce => \N__41096\,
            sr => \N__48622\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41099\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49025\,
            ce => \N__41096\,
            sr => \N__48622\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48072\,
            in1 => \N__48221\,
            in2 => \_gnd_net_\,
            in3 => \N__49568\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49020\,
            ce => \N__48718\,
            sr => \N__48628\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49567\,
            in1 => \N__41007\,
            in2 => \_gnd_net_\,
            in3 => \N__40991\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49020\,
            ce => \N__48718\,
            sr => \N__48628\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43616\,
            in1 => \N__43895\,
            in2 => \_gnd_net_\,
            in3 => \N__49570\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49020\,
            ce => \N__48718\,
            sr => \N__48628\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40919\,
            in1 => \N__43866\,
            in2 => \_gnd_net_\,
            in3 => \N__49571\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49020\,
            ce => \N__48718\,
            sr => \N__48628\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43585\,
            in1 => \N__43554\,
            in2 => \_gnd_net_\,
            in3 => \N__49569\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49020\,
            ce => \N__48718\,
            sr => \N__48628\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47631\,
            in1 => \N__47890\,
            in2 => \_gnd_net_\,
            in3 => \N__49554\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49016\,
            ce => \N__48716\,
            sr => \N__48635\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41425\,
            in1 => \N__44704\,
            in2 => \N__42476\,
            in3 => \N__45622\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45621\,
            in1 => \N__41855\,
            in2 => \_gnd_net_\,
            in3 => \N__41424\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41853\,
            in1 => \N__44298\,
            in2 => \_gnd_net_\,
            in3 => \N__41400\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__41852\,
            in1 => \N__41379\,
            in2 => \_gnd_net_\,
            in3 => \N__41363\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45687\,
            in1 => \N__41854\,
            in2 => \_gnd_net_\,
            in3 => \N__41325\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41856\,
            in1 => \N__45549\,
            in2 => \_gnd_net_\,
            in3 => \N__41301\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41285\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46245\,
            in1 => \N__41861\,
            in2 => \_gnd_net_\,
            in3 => \N__41199\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__41857\,
            in1 => \N__41181\,
            in2 => \_gnd_net_\,
            in3 => \N__44356\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46176\,
            in1 => \N__41862\,
            in2 => \_gnd_net_\,
            in3 => \N__41160\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41860\,
            in1 => \N__45151\,
            in2 => \_gnd_net_\,
            in3 => \N__41565\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45548\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__41858\,
            in1 => \_gnd_net_\,
            in2 => \N__44223\,
            in3 => \N__41532\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41508\,
            in1 => \N__41859\,
            in2 => \_gnd_net_\,
            in3 => \N__44137\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45231\,
            in1 => \N__41844\,
            in2 => \_gnd_net_\,
            in3 => \N__41490\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44355\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46854\,
            in1 => \N__41846\,
            in2 => \_gnd_net_\,
            in3 => \N__41460\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44288\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41843\,
            in1 => \N__45393\,
            in2 => \_gnd_net_\,
            in3 => \N__41748\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45819\,
            in1 => \N__41845\,
            in2 => \_gnd_net_\,
            in3 => \N__41727\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44136\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44725\,
            in1 => \N__46641\,
            in2 => \_gnd_net_\,
            in3 => \N__41694\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__41803\,
            in1 => \N__41676\,
            in2 => \_gnd_net_\,
            in3 => \N__46035\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__45963\,
            in1 => \N__41646\,
            in2 => \_gnd_net_\,
            in3 => \N__41804\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46782\,
            in1 => \N__41806\,
            in2 => \_gnd_net_\,
            in3 => \N__41622\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46497\,
            in1 => \N__44726\,
            in2 => \_gnd_net_\,
            in3 => \N__41598\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46101\,
            in1 => \N__41802\,
            in2 => \_gnd_net_\,
            in3 => \N__42570\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__41805\,
            in1 => \_gnd_net_\,
            in2 => \N__45891\,
            in3 => \N__42546\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__46408\,
            in1 => \N__44756\,
            in2 => \N__42515\,
            in3 => \N__42399\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44753\,
            in1 => \N__46407\,
            in2 => \_gnd_net_\,
            in3 => \N__42510\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44757\,
            in2 => \_gnd_net_\,
            in3 => \N__42398\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44754\,
            in1 => \N__45748\,
            in2 => \N__42465\,
            in3 => \N__41878\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__45749\,
            in1 => \N__44755\,
            in2 => \N__41879\,
            in3 => \N__42403\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__41807\,
            in1 => \N__45747\,
            in2 => \_gnd_net_\,
            in3 => \N__41874\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47121\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49117\,
            ce => \N__47164\,
            sr => \N__48523\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45945\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45375\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46228\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45873\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45294\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45221\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46772\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46158\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46302\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46836\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46478\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45800\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45739\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46697\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46623\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42758\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47207\,
            in2 => \N__42689\,
            in3 => \N__43083\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47738\,
            in2 => \N__42680\,
            in3 => \N__43058\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42947\,
            in2 => \N__42941\,
            in3 => \N__43033\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42932\,
            in2 => \N__42926\,
            in3 => \N__43313\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42917\,
            in2 => \N__47336\,
            in3 => \N__43295\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43277\,
            in1 => \N__47018\,
            in2 => \N__42911\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42902\,
            in2 => \N__42896\,
            in3 => \N__43259\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42884\,
            in2 => \N__42872\,
            in3 => \N__43241\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42860\,
            in2 => \N__42848\,
            in3 => \N__43223\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42839\,
            in2 => \N__42827\,
            in3 => \N__43205\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43013\,
            in2 => \N__43001\,
            in3 => \N__43184\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42992\,
            in2 => \N__42980\,
            in3 => \N__43403\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43820\,
            in2 => \N__42971\,
            in3 => \N__43385\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43367\,
            in1 => \N__46892\,
            in2 => \N__42962\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42953\,
            in2 => \N__47615\,
            in3 => \N__43349\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47012\,
            in2 => \N__46925\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47510\,
            in2 => \N__47558\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47318\,
            in2 => \N__47270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43166\,
            in2 => \N__43154\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47402\,
            in2 => \N__47462\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48191\,
            in2 => \N__47975\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43625\,
            in2 => \N__43676\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43139\,
            in2 => \N__43133\,
            in3 => \N__43109\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43106\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43090\,
            in2 => \N__43067\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49998\,
            in1 => \N__43057\,
            in2 => \_gnd_net_\,
            in3 => \N__43043\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__49975\,
            in1 => \N__43040\,
            in2 => \N__43034\,
            in3 => \N__43016\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49999\,
            in1 => \N__43312\,
            in2 => \_gnd_net_\,
            in3 => \N__43298\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49976\,
            in1 => \N__43294\,
            in2 => \_gnd_net_\,
            in3 => \N__43280\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50000\,
            in1 => \N__43276\,
            in2 => \_gnd_net_\,
            in3 => \N__43262\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49977\,
            in1 => \N__43258\,
            in2 => \_gnd_net_\,
            in3 => \N__43244\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50001\,
            in1 => \N__43240\,
            in2 => \_gnd_net_\,
            in3 => \N__43226\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49063\,
            ce => 'H',
            sr => \N__48568\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49981\,
            in1 => \N__43222\,
            in2 => \_gnd_net_\,
            in3 => \N__43208\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49961\,
            in1 => \N__43201\,
            in2 => \_gnd_net_\,
            in3 => \N__43187\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49978\,
            in1 => \N__43183\,
            in2 => \_gnd_net_\,
            in3 => \N__43169\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49962\,
            in1 => \N__43402\,
            in2 => \_gnd_net_\,
            in3 => \N__43388\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49979\,
            in1 => \N__43384\,
            in2 => \_gnd_net_\,
            in3 => \N__43370\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49963\,
            in1 => \N__43366\,
            in2 => \_gnd_net_\,
            in3 => \N__43352\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49980\,
            in1 => \N__43345\,
            in2 => \_gnd_net_\,
            in3 => \N__43331\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49964\,
            in1 => \N__46948\,
            in2 => \_gnd_net_\,
            in3 => \N__43328\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49057\,
            ce => 'H',
            sr => \N__48579\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49953\,
            in1 => \N__46975\,
            in2 => \_gnd_net_\,
            in3 => \N__43325\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50048\,
            in1 => \N__47543\,
            in2 => \_gnd_net_\,
            in3 => \N__43322\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49954\,
            in1 => \N__47527\,
            in2 => \_gnd_net_\,
            in3 => \N__43319\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50049\,
            in1 => \N__47310\,
            in2 => \_gnd_net_\,
            in3 => \N__43316\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49955\,
            in1 => \N__47286\,
            in2 => \_gnd_net_\,
            in3 => \N__43466\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50050\,
            in1 => \N__43462\,
            in2 => \_gnd_net_\,
            in3 => \N__43445\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49956\,
            in1 => \N__43441\,
            in2 => \_gnd_net_\,
            in3 => \N__43424\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50051\,
            in1 => \N__47418\,
            in2 => \_gnd_net_\,
            in3 => \N__43421\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49050\,
            ce => 'H',
            sr => \N__48587\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49957\,
            in1 => \N__47445\,
            in2 => \_gnd_net_\,
            in3 => \N__43418\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50053\,
            in1 => \N__48005\,
            in2 => \_gnd_net_\,
            in3 => \N__43415\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49958\,
            in1 => \N__47990\,
            in2 => \_gnd_net_\,
            in3 => \N__43412\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50054\,
            in1 => \N__43661\,
            in2 => \_gnd_net_\,
            in3 => \N__43409\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49959\,
            in1 => \N__43641\,
            in2 => \_gnd_net_\,
            in3 => \N__43406\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50055\,
            in1 => \N__43727\,
            in2 => \_gnd_net_\,
            in3 => \N__43709\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49960\,
            in1 => \N__43690\,
            in2 => \_gnd_net_\,
            in3 => \N__43706\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49043\,
            ce => 'H',
            sr => \N__48595\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__43659\,
            in1 => \N__43642\,
            in2 => \N__43598\,
            in3 => \N__43538\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__43537\,
            in1 => \N__43660\,
            in2 => \N__43646\,
            in3 => \N__43594\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43893\,
            in1 => \N__43612\,
            in2 => \_gnd_net_\,
            in3 => \N__49454\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49456\,
            in1 => \_gnd_net_\,
            in2 => \N__43601\,
            in3 => \N__43894\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49035\,
            ce => \N__50032\,
            sr => \N__48605\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49455\,
            in1 => \N__43586\,
            in2 => \_gnd_net_\,
            in3 => \N__43562\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49035\,
            ce => \N__50032\,
            sr => \N__48605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43515\,
            in1 => \N__43482\,
            in2 => \N__47678\,
            in3 => \N__47356\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43892\,
            in1 => \N__50162\,
            in2 => \N__47948\,
            in3 => \N__43862\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43841\,
            in1 => \N__49616\,
            in2 => \_gnd_net_\,
            in3 => \N__47808\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49030\,
            ce => \N__50033\,
            sr => \N__48614\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49637\,
            in1 => \N__48143\,
            in2 => \_gnd_net_\,
            in3 => \N__47493\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47635\,
            in1 => \N__47886\,
            in2 => \_gnd_net_\,
            in3 => \N__49636\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49638\,
            in1 => \N__50259\,
            in2 => \_gnd_net_\,
            in3 => \N__50235\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49635\,
            in1 => \N__47094\,
            in2 => \_gnd_net_\,
            in3 => \N__47040\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43808\,
            in2 => \N__43772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_7_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45075\,
            in2 => \N__43751\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43742\,
            in2 => \N__45096\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45079\,
            in2 => \N__43976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43967\,
            in2 => \N__45097\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45083\,
            in2 => \N__43961\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43952\,
            in2 => \N__45098\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45087\,
            in2 => \N__43946\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44965\,
            in2 => \N__43937\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43928\,
            in2 => \N__45039\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44953\,
            in2 => \N__43913\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43904\,
            in2 => \N__45036\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44957\,
            in2 => \N__44036\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44027\,
            in2 => \N__45037\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44961\,
            in2 => \N__44021\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44012\,
            in2 => \N__45038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45059\,
            in2 => \N__44006\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43997\,
            in2 => \N__45092\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45063\,
            in2 => \N__43991\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43982\,
            in2 => \N__45093\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45067\,
            in2 => \N__44111\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44102\,
            in2 => \N__45094\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45071\,
            in2 => \N__44093\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44084\,
            in2 => \N__45095\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45046\,
            in2 => \N__44078\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44063\,
            in2 => \N__45089\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45050\,
            in2 => \N__44057\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44042\,
            in2 => \N__45090\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45054\,
            in2 => \N__45119\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45107\,
            in2 => \N__45091\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45058\,
            in2 => \N__44774\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44727\,
            in2 => \_gnd_net_\,
            in3 => \N__44474\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44392\,
            in2 => \N__44260\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44336\,
            in2 => \N__44182\,
            in3 => \N__44264\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45721\,
            in2 => \N__44261\,
            in3 => \N__44186\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45646\,
            in2 => \N__44183\,
            in3 => \N__44114\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45583\,
            in2 => \N__45725\,
            in3 => \N__45650\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45647\,
            in2 => \N__45505\,
            in3 => \N__45587\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45584\,
            in2 => \N__45439\,
            in3 => \N__45509\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45352\,
            in2 => \N__45506\,
            in3 => \N__45443\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__49124\,
            ce => \N__47167\,
            sr => \N__48520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45271\,
            in2 => \N__45440\,
            in3 => \N__45359\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45193\,
            in2 => \N__45356\,
            in3 => \N__45278\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46279\,
            in2 => \N__45275\,
            in3 => \N__45200\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46213\,
            in2 => \N__45197\,
            in3 => \N__45122\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46135\,
            in2 => \N__46283\,
            in3 => \N__46217\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46214\,
            in2 => \N__46063\,
            in3 => \N__46142\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45994\,
            in2 => \N__46139\,
            in3 => \N__46067\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45919\,
            in2 => \N__46064\,
            in3 => \N__46004\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__49118\,
            ce => \N__47165\,
            sr => \N__48524\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45850\,
            in2 => \N__46001\,
            in3 => \N__45929\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45772\,
            in2 => \N__45926\,
            in3 => \N__45857\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46885\,
            in2 => \N__45854\,
            in3 => \N__45779\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46816\,
            in2 => \N__45776\,
            in3 => \N__45728\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46886\,
            in2 => \N__46750\,
            in3 => \N__46820\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46817\,
            in2 => \N__46672\,
            in3 => \N__46754\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46597\,
            in2 => \N__46751\,
            in3 => \N__46676\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46528\,
            in2 => \N__46673\,
            in3 => \N__46607\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__49108\,
            ce => \N__47162\,
            sr => \N__48526\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46432\,
            in2 => \N__46604\,
            in3 => \N__46538\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__49101\,
            ce => \N__47161\,
            sr => \N__48530\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46351\,
            in2 => \N__46535\,
            in3 => \N__46457\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__49101\,
            ce => \N__47161\,
            sr => \N__48530\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46454\,
            in2 => \N__46436\,
            in3 => \N__46376\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__49101\,
            ce => \N__47161\,
            sr => \N__48530\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46373\,
            in2 => \N__46355\,
            in3 => \N__46286\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__49101\,
            ce => \N__47161\,
            sr => \N__48530\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47138\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47096\,
            in1 => \N__47048\,
            in2 => \_gnd_net_\,
            in3 => \N__49640\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49093\,
            ce => \N__50066\,
            sr => \N__48536\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__46982\,
            in1 => \N__47570\,
            in2 => \N__46961\,
            in3 => \N__46934\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49584\,
            in1 => \N__48178\,
            in2 => \_gnd_net_\,
            in3 => \N__46996\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__48179\,
            in1 => \_gnd_net_\,
            in2 => \N__46985\,
            in3 => \N__49587\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49084\,
            ce => \N__50034\,
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__46981\,
            in1 => \N__47569\,
            in2 => \N__46960\,
            in3 => \N__46933\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47851\,
            in1 => \N__49585\,
            in2 => \_gnd_net_\,
            in3 => \N__46906\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49586\,
            in1 => \_gnd_net_\,
            in2 => \N__46895\,
            in3 => \N__47852\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49084\,
            ce => \N__50034\,
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__47425\,
            in1 => \N__47453\,
            in2 => \N__47726\,
            in3 => \N__47345\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__47344\,
            in1 => \N__47452\,
            in2 => \N__47429\,
            in3 => \N__47722\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47376\,
            in1 => \N__47392\,
            in2 => \_gnd_net_\,
            in3 => \N__49629\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49630\,
            in1 => \_gnd_net_\,
            in2 => \N__47381\,
            in3 => \N__47377\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49076\,
            ce => \N__50062\,
            sr => \N__48549\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49714\,
            in1 => \N__49666\,
            in2 => \_gnd_net_\,
            in3 => \N__49631\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49076\,
            ce => \N__50062\,
            sr => \N__48549\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__47579\,
            in1 => \N__47312\,
            in2 => \N__47294\,
            in3 => \N__47648\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__47578\,
            in1 => \N__47311\,
            in2 => \N__47293\,
            in3 => \N__47647\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47258\,
            in1 => \N__47234\,
            in2 => \_gnd_net_\,
            in3 => \N__49619\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49069\,
            ce => \N__49990\,
            sr => \N__48557\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49618\,
            in1 => \N__47195\,
            in2 => \_gnd_net_\,
            in3 => \N__47768\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49069\,
            ce => \N__49990\,
            sr => \N__48557\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47914\,
            in1 => \N__47960\,
            in2 => \_gnd_net_\,
            in3 => \N__49592\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49064\,
            ce => \N__50005\,
            sr => \N__48569\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47711\,
            in1 => \N__47687\,
            in2 => \_gnd_net_\,
            in3 => \N__49591\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49064\,
            ce => \N__50005\,
            sr => \N__48569\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47639\,
            in1 => \N__47891\,
            in2 => \_gnd_net_\,
            in3 => \N__49589\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49064\,
            ce => \N__50005\,
            sr => \N__48569\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49588\,
            in1 => \N__47603\,
            in2 => \_gnd_net_\,
            in3 => \N__48111\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49064\,
            ce => \N__50005\,
            sr => \N__48569\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49741\,
            in1 => \N__49778\,
            in2 => \_gnd_net_\,
            in3 => \N__49590\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49064\,
            ce => \N__50005\,
            sr => \N__48569\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__47541\,
            in1 => \N__47523\,
            in2 => \N__47474\,
            in3 => \N__48200\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__48199\,
            in1 => \N__47542\,
            in2 => \N__47528\,
            in3 => \N__47470\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49615\,
            in1 => \N__47500\,
            in2 => \_gnd_net_\,
            in3 => \N__48148\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49058\,
            ce => \N__50047\,
            sr => \N__48580\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48073\,
            in1 => \N__48214\,
            in2 => \_gnd_net_\,
            in3 => \N__49613\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49614\,
            in1 => \_gnd_net_\,
            in2 => \N__48203\,
            in3 => \N__48074\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49058\,
            ce => \N__50047\,
            sr => \N__48580\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__50144\,
            in1 => \N__48004\,
            in2 => \N__50213\,
            in3 => \N__47989\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48168\,
            in1 => \N__48147\,
            in2 => \N__48113\,
            in3 => \N__48066\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48044\,
            in1 => \N__48035\,
            in2 => \N__48026\,
            in3 => \N__47774\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__50143\,
            in1 => \N__48003\,
            in2 => \N__50212\,
            in3 => \N__47988\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47913\,
            in1 => \N__47958\,
            in2 => \_gnd_net_\,
            in3 => \N__49593\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47885\,
            in1 => \N__47844\,
            in2 => \N__49777\,
            in3 => \N__47801\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50267\,
            in1 => \N__50237\,
            in2 => \_gnd_net_\,
            in3 => \N__49458\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49044\,
            ce => \N__49983\,
            sr => \N__48596\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50198\,
            in1 => \N__50173\,
            in2 => \_gnd_net_\,
            in3 => \N__49457\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49044\,
            ce => \N__49983\,
            sr => \N__48596\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50135\,
            in2 => \_gnd_net_\,
            in3 => \N__50100\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49659\,
            in1 => \N__49713\,
            in2 => \_gnd_net_\,
            in3 => \N__49617\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49734\,
            in1 => \N__49773\,
            in2 => \_gnd_net_\,
            in3 => \N__49639\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49715\,
            in1 => \N__49667\,
            in2 => \_gnd_net_\,
            in3 => \N__49555\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49045\,
            ce => \N__48721\,
            sr => \N__48615\
        );
end \INTERFACE\;
